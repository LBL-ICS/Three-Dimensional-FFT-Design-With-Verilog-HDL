module cmplx_adj(
  input  [31:0] io_in_Re,
  input  [31:0] io_in_Im,
  input  [7:0]  io_in_adj,
  input         io_is_neg,
  input         io_is_flip,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  wire  sign_0 = io_in_Re[31]; // @[FFTDesigns.scala 4716:24]
  wire  sign_1 = io_in_Im[31]; // @[FFTDesigns.scala 4717:24]
  wire [7:0] exp_0 = io_in_Re[30:23]; // @[FFTDesigns.scala 4719:23]
  wire [7:0] exp_1 = io_in_Im[30:23]; // @[FFTDesigns.scala 4720:23]
  wire [22:0] frac_0 = io_in_Re[22:0]; // @[FFTDesigns.scala 4722:24]
  wire [22:0] frac_1 = io_in_Im[22:0]; // @[FFTDesigns.scala 4723:24]
  wire  new_sign_0 = io_is_neg ? ~sign_0 : sign_0; // @[FFTDesigns.scala 4725:20 4726:19 4729:19]
  wire  new_sign_1 = io_is_neg ? ~sign_1 : sign_1; // @[FFTDesigns.scala 4725:20 4727:19 4730:19]
  wire [7:0] _new_exp_0_T_1 = exp_0 - io_in_adj; // @[FFTDesigns.scala 4734:28]
  wire [7:0] new_exp_0 = exp_0 != 8'h0 ? _new_exp_0_T_1 : exp_0; // @[FFTDesigns.scala 4733:25 4734:18 4736:18]
  wire [7:0] _new_exp_1_T_1 = exp_1 - io_in_adj; // @[FFTDesigns.scala 4739:28]
  wire [7:0] new_exp_1 = exp_1 != 8'h0 ? _new_exp_1_T_1 : exp_1; // @[FFTDesigns.scala 4738:26 4739:18 4741:18]
  wire  _io_out_Re_T = ~new_sign_1; // @[FFTDesigns.scala 4745:21]
  wire [31:0] _io_out_Re_T_2 = {_io_out_Re_T,new_exp_1,frac_1}; // @[FFTDesigns.scala 4745:49]
  wire [31:0] _io_out_Im_T_1 = {new_sign_0,new_exp_0,frac_0}; // @[FFTDesigns.scala 4746:48]
  wire [31:0] _io_out_Im_T_3 = {new_sign_1,new_exp_1,frac_1}; // @[FFTDesigns.scala 4749:48]
  assign io_out_Re = io_is_flip ? _io_out_Re_T_2 : _io_out_Im_T_1; // @[FFTDesigns.scala 4744:21 4745:17 4748:17]
  assign io_out_Im = io_is_flip ? _io_out_Im_T_1 : _io_out_Im_T_3; // @[FFTDesigns.scala 4744:21 4746:17 4749:17]
endmodule
module full_subber(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[Arithmetic.scala 72:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[Arithmetic.scala 72:34]
  wire [8:0] result = _result_T_2[8:0]; // @[Arithmetic.scala 71:22 72:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 73:23]
  assign io_out_c = result[8]; // @[Arithmetic.scala 74:23]
endmodule
module twoscomplement(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _x_T = ~io_in; // @[Arithmetic.scala 28:16]
  assign io_out = 8'h1 + _x_T; // @[Arithmetic.scala 28:14]
endmodule
module full_adder(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 58:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 58:34]
  wire [24:0] result = _result_T_1[24:0]; // @[Arithmetic.scala 57:22 58:12]
  assign io_out_s = result[23:0]; // @[Arithmetic.scala 59:23]
  assign io_out_c = result[24]; // @[Arithmetic.scala 60:23]
endmodule
module twoscomplement_1(
  input  [23:0] io_in,
  output [23:0] io_out
);
  wire [23:0] _x_T = ~io_in; // @[Arithmetic.scala 28:16]
  assign io_out = 24'h1 + _x_T; // @[Arithmetic.scala 28:14]
endmodule
module shifter(
  input  [23:0] io_in_a,
  input  [4:0]  io_in_b,
  output [23:0] io_out_s
);
  wire [23:0] _result_T = io_in_a >> io_in_b; // @[Arithmetic.scala 42:25]
  wire [54:0] _GEN_0 = {{31'd0}, _result_T}; // @[Arithmetic.scala 41:26 42:14 44:14]
  assign io_out_s = _GEN_0[23:0]; // @[Arithmetic.scala 39:22]
endmodule
module leadingOneDetector(
  input  [23:0] io_in,
  output [4:0]  io_out
);
  wire [1:0] _hotValue_T = io_in[1] ? 2'h2 : 2'h1; // @[Mux.scala 47:70]
  wire [1:0] _hotValue_T_1 = io_in[2] ? 2'h3 : _hotValue_T; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_2 = io_in[3] ? 3'h4 : {{1'd0}, _hotValue_T_1}; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_3 = io_in[4] ? 3'h5 : _hotValue_T_2; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_4 = io_in[5] ? 3'h6 : _hotValue_T_3; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_5 = io_in[6] ? 3'h7 : _hotValue_T_4; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_6 = io_in[7] ? 4'h8 : {{1'd0}, _hotValue_T_5}; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_7 = io_in[8] ? 4'h9 : _hotValue_T_6; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_8 = io_in[9] ? 4'ha : _hotValue_T_7; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_9 = io_in[10] ? 4'hb : _hotValue_T_8; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_10 = io_in[11] ? 4'hc : _hotValue_T_9; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_11 = io_in[12] ? 4'hd : _hotValue_T_10; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_12 = io_in[13] ? 4'he : _hotValue_T_11; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_13 = io_in[14] ? 4'hf : _hotValue_T_12; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_14 = io_in[15] ? 5'h10 : {{1'd0}, _hotValue_T_13}; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_15 = io_in[16] ? 5'h11 : _hotValue_T_14; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_16 = io_in[17] ? 5'h12 : _hotValue_T_15; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_17 = io_in[18] ? 5'h13 : _hotValue_T_16; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_18 = io_in[19] ? 5'h14 : _hotValue_T_17; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_19 = io_in[20] ? 5'h15 : _hotValue_T_18; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_20 = io_in[21] ? 5'h16 : _hotValue_T_19; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_21 = io_in[22] ? 5'h17 : _hotValue_T_20; // @[Mux.scala 47:70]
  assign io_out = io_in[23] ? 5'h18 : _hotValue_T_21; // @[Mux.scala 47:70]
endmodule
module FP_adder(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 76:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 76:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 76:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 76:24]
  wire [7:0] complement_io_in; // @[FPArithmetic.scala 82:28]
  wire [7:0] complement_io_out; // @[FPArithmetic.scala 82:28]
  wire [23:0] adder_io_in_a; // @[FPArithmetic.scala 86:23]
  wire [23:0] adder_io_in_b; // @[FPArithmetic.scala 86:23]
  wire [23:0] adder_io_out_s; // @[FPArithmetic.scala 86:23]
  wire  adder_io_out_c; // @[FPArithmetic.scala 86:23]
  wire [23:0] complementN_0_io_in; // @[FPArithmetic.scala 92:31]
  wire [23:0] complementN_0_io_out; // @[FPArithmetic.scala 92:31]
  wire [23:0] complementN_1_io_in; // @[FPArithmetic.scala 94:31]
  wire [23:0] complementN_1_io_out; // @[FPArithmetic.scala 94:31]
  wire [23:0] shifter_io_in_a; // @[FPArithmetic.scala 98:25]
  wire [4:0] shifter_io_in_b; // @[FPArithmetic.scala 98:25]
  wire [23:0] shifter_io_out_s; // @[FPArithmetic.scala 98:25]
  wire [23:0] complementN_2_io_in; // @[FPArithmetic.scala 143:31]
  wire [23:0] complementN_2_io_out; // @[FPArithmetic.scala 143:31]
  wire [23:0] leadingOneFinder_io_in; // @[FPArithmetic.scala 163:34]
  wire [4:0] leadingOneFinder_io_out; // @[FPArithmetic.scala 163:34]
  wire [7:0] subber2_io_in_a; // @[FPArithmetic.scala 165:25]
  wire [7:0] subber2_io_in_b; // @[FPArithmetic.scala 165:25]
  wire [7:0] subber2_io_out_s; // @[FPArithmetic.scala 165:25]
  wire  subber2_io_out_c; // @[FPArithmetic.scala 165:25]
  wire  sign_0 = io_in_a[31]; // @[FPArithmetic.scala 38:23]
  wire  sign_1 = io_in_b[31]; // @[FPArithmetic.scala 39:23]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 43:62]
  wire [8:0] _GEN_31 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 43:34]
  wire [8:0] _GEN_0 = _GEN_31 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 43:68 44:14 46:14]
  wire [8:0] _GEN_32 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 48:34]
  wire [8:0] _GEN_1 = _GEN_32 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 48:68 49:14 51:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 56:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 57:23]
  wire [23:0] whole_frac_0 = {1'h1,frac_0}; // @[FPArithmetic.scala 61:26]
  wire [23:0] whole_frac_1 = {1'h1,frac_1}; // @[FPArithmetic.scala 62:26]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 42:19]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 42:19]
  wire [7:0] out_exp = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 104:34 105:15 115:15]
  wire [7:0] sub_exp = subber_io_out_c ? complement_io_out : subber_io_out_s; // @[FPArithmetic.scala 104:34 106:15 116:15]
  wire  out_s = subber_io_out_c ? sign_1 : sign_0; // @[FPArithmetic.scala 104:34 107:13 117:13]
  wire [22:0] out_frac = subber_io_out_c ? frac_1 : frac_0; // @[FPArithmetic.scala 104:34 108:16 118:16]
  wire [23:0] _GEN_8 = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 104:34 112:21 87:19]
  wire [23:0] _GEN_9 = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 104:34 88:19 122:21]
  wire  _new_s_T = ~adder_io_out_c; // @[FPArithmetic.scala 138:15]
  wire  _D_T_1 = sign_0 ^ sign_1; // @[FPArithmetic.scala 151:39]
  wire  D = _new_s_T | sign_0 ^ sign_1; // @[FPArithmetic.scala 151:28]
  wire  E = _new_s_T & ~adder_io_out_s[23] | _new_s_T & ~_D_T_1 | adder_io_out_c & adder_io_out_s[23] & _D_T_1; // @[FPArithmetic.scala 154:99]
  wire  _GEN_25 = sub_exp >= 8'h17 ? out_s : ~adder_io_out_c & sign_0 | sign_0 & sign_1 | ~adder_io_out_c & sign_1; // @[FPArithmetic.scala 138:11 173:39 174:13]
  wire  new_s = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 1'h0 : _GEN_25; // @[FPArithmetic.scala 169:62 170:13]
  wire [23:0] adder_result = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 157:18 158:47 159:20]
  wire [4:0] _subber2_io_in_b_T_1 = 5'h18 - leadingOneFinder_io_out; // @[FPArithmetic.scala 167:42]
  wire [8:0] _GEN_33 = {{1'd0}, out_exp}; // @[FPArithmetic.scala 181:20]
  wire [23:0] _new_out_frac_T_2 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 183:51]
  wire [7:0] _new_out_exp_T_3 = out_exp + 8'h1; // @[FPArithmetic.scala 185:32]
  wire [8:0] _GEN_13 = _GEN_33 == _T_2 ? _T_2 : {{1'd0}, _new_out_exp_T_3}; // @[FPArithmetic.scala 181:56 182:21 185:21]
  wire [23:0] _GEN_14 = _GEN_33 == _T_2 ? _new_out_frac_T_2 : {{1'd0}, adder_result[23:1]}; // @[FPArithmetic.scala 181:56 183:22 186:22]
  wire [53:0] _GEN_2 = {{31'd0}, adder_result[22:0]}; // @[FPArithmetic.scala 197:57]
  wire [53:0] _new_out_frac_T_7 = _GEN_2 << _subber2_io_in_b_T_1; // @[FPArithmetic.scala 197:57]
  wire [7:0] _GEN_15 = subber2_io_out_c ? 8'h1 : subber2_io_out_s; // @[FPArithmetic.scala 192:39 193:23 196:23]
  wire [53:0] _GEN_16 = subber2_io_out_c ? 54'h400000 : _new_out_frac_T_7; // @[FPArithmetic.scala 192:39 194:24 197:24]
  wire [7:0] _GEN_17 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:0
    ]) ? 8'h0 : _GEN_15; // @[FPArithmetic.scala 189:141 190:21]
  wire [53:0] _GEN_18 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:
    0]) ? 54'h0 : _GEN_16; // @[FPArithmetic.scala 189:141 139:18]
  wire [7:0] _GEN_19 = D ? _GEN_17 : 8'h0; // @[FPArithmetic.scala 140:17 188:26]
  wire [53:0] _GEN_20 = D ? _GEN_18 : 54'h0; // @[FPArithmetic.scala 139:18 188:26]
  wire [8:0] _GEN_21 = ~D ? _GEN_13 : {{1'd0}, _GEN_19}; // @[FPArithmetic.scala 180:26]
  wire [53:0] _GEN_22 = ~D ? {{30'd0}, _GEN_14} : _GEN_20; // @[FPArithmetic.scala 180:26]
  wire [8:0] _GEN_23 = E ? {{1'd0}, out_exp} : _GEN_21; // @[FPArithmetic.scala 177:26 178:19]
  wire [53:0] _GEN_24 = E ? {{31'd0}, adder_result[22:0]} : _GEN_22; // @[FPArithmetic.scala 177:26 179:20]
  wire [53:0] _GEN_26 = sub_exp >= 8'h17 ? {{31'd0}, out_frac} : _GEN_24; // @[FPArithmetic.scala 173:39 175:20]
  wire [8:0] _GEN_27 = sub_exp >= 8'h17 ? {{1'd0}, out_exp} : _GEN_23; // @[FPArithmetic.scala 173:39 176:19]
  wire [8:0] _GEN_29 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 9'h0 : _GEN_27; // @[FPArithmetic.scala 169:62 171:19]
  wire [53:0] _GEN_30 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 54'h0 : _GEN_26; // @[FPArithmetic.scala 169:62 172:20]
  reg [31:0] reg_out_s; // @[FPArithmetic.scala 201:28]
  wire [7:0] new_out_exp = _GEN_29[7:0]; // @[FPArithmetic.scala 137:27]
  wire [22:0] new_out_frac = _GEN_30[22:0]; // @[FPArithmetic.scala 136:28]
  wire [31:0] _reg_out_s_T_1 = {new_s,new_out_exp,new_out_frac}; // @[FPArithmetic.scala 203:39]
  full_subber subber ( // @[FPArithmetic.scala 76:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complement ( // @[FPArithmetic.scala 82:28]
    .io_in(complement_io_in),
    .io_out(complement_io_out)
  );
  full_adder adder ( // @[FPArithmetic.scala 86:23]
    .io_in_a(adder_io_in_a),
    .io_in_b(adder_io_in_b),
    .io_out_s(adder_io_out_s),
    .io_out_c(adder_io_out_c)
  );
  twoscomplement_1 complementN_0 ( // @[FPArithmetic.scala 92:31]
    .io_in(complementN_0_io_in),
    .io_out(complementN_0_io_out)
  );
  twoscomplement_1 complementN_1 ( // @[FPArithmetic.scala 94:31]
    .io_in(complementN_1_io_in),
    .io_out(complementN_1_io_out)
  );
  shifter shifter ( // @[FPArithmetic.scala 98:25]
    .io_in_a(shifter_io_in_a),
    .io_in_b(shifter_io_in_b),
    .io_out_s(shifter_io_out_s)
  );
  twoscomplement_1 complementN_2 ( // @[FPArithmetic.scala 143:31]
    .io_in(complementN_2_io_in),
    .io_out(complementN_2_io_out)
  );
  leadingOneDetector leadingOneFinder ( // @[FPArithmetic.scala 163:34]
    .io_in(leadingOneFinder_io_in),
    .io_out(leadingOneFinder_io_out)
  );
  full_subber subber2 ( // @[FPArithmetic.scala 165:25]
    .io_in_a(subber2_io_in_a),
    .io_in_b(subber2_io_in_b),
    .io_out_s(subber2_io_out_s),
    .io_out_c(subber2_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FPArithmetic.scala 205:14]
  assign subber_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 42:19]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 42:19]
  assign complement_io_in = subber_io_out_s; // @[FPArithmetic.scala 83:22]
  assign adder_io_in_a = sign_0 & ~sign_1 ? complementN_0_io_out : _GEN_8; // @[FPArithmetic.scala 127:45 128:21]
  assign adder_io_in_b = sign_1 & ~sign_0 ? complementN_1_io_out : _GEN_9; // @[FPArithmetic.scala 131:45 132:21]
  assign complementN_0_io_in = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 104:34 112:21 87:19]
  assign complementN_1_io_in = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 104:34 88:19 122:21]
  assign shifter_io_in_a = subber_io_out_c ? whole_frac_0 : whole_frac_1; // @[FPArithmetic.scala 104:34 109:23 119:23]
  assign shifter_io_in_b = sub_exp[4:0];
  assign complementN_2_io_in = adder_io_out_s; // @[FPArithmetic.scala 144:25]
  assign leadingOneFinder_io_in = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 157:18 158:47 159:20]
  assign subber2_io_in_a = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 104:34 105:15 115:15]
  assign subber2_io_in_b = {{3'd0}, _subber2_io_in_b_T_1}; // @[FPArithmetic.scala 167:21]
  always @(posedge clock) begin
    if (reset) begin // @[FPArithmetic.scala 201:28]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 201:28]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FPArithmetic.scala 203:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_out_s = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexAdder(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_adder_clock; // @[FPComplex.scala 21:25]
  wire  FP_adder_reset; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 21:25]
  wire  FP_adder_1_clock; // @[FPComplex.scala 21:25]
  wire  FP_adder_1_reset; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_in_a; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_in_b; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_out_s; // @[FPComplex.scala 21:25]
  FP_adder FP_adder ( // @[FPComplex.scala 21:25]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_adder FP_adder_1 ( // @[FPComplex.scala 21:25]
    .clock(FP_adder_1_clock),
    .reset(FP_adder_1_reset),
    .io_in_a(FP_adder_1_io_in_a),
    .io_in_b(FP_adder_1_io_in_b),
    .io_out_s(FP_adder_1_io_out_s)
  );
  assign io_out_s_Re = FP_adder_io_out_s; // @[FPComplex.scala 28:17]
  assign io_out_s_Im = FP_adder_1_io_out_s; // @[FPComplex.scala 29:17]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = io_in_a_Re; // @[FPComplex.scala 24:23]
  assign FP_adder_io_in_b = io_in_b_Re; // @[FPComplex.scala 25:23]
  assign FP_adder_1_clock = clock;
  assign FP_adder_1_reset = reset;
  assign FP_adder_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 26:23]
  assign FP_adder_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 27:23]
endmodule
module FPComplexMultiAdder(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  wire  FPComplexAdder_clock; // @[FPComplex.scala 524:30]
  wire  FPComplexAdder_reset; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_in_a_Re; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_in_a_Im; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_in_b_Re; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_in_b_Im; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_out_s_Re; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_out_s_Im; // @[FPComplex.scala 524:30]
  FPComplexAdder FPComplexAdder ( // @[FPComplex.scala 524:30]
    .clock(FPComplexAdder_clock),
    .reset(FPComplexAdder_reset),
    .io_in_a_Re(FPComplexAdder_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_io_out_s_Im)
  );
  assign io_out_Re = FPComplexAdder_io_out_s_Re; // @[FPComplex.scala 642:16]
  assign io_out_Im = FPComplexAdder_io_out_s_Im; // @[FPComplex.scala 642:16]
  assign FPComplexAdder_clock = clock;
  assign FPComplexAdder_reset = reset;
  assign FPComplexAdder_io_in_a_Re = io_in_0_Re; // @[FPComplex.scala 604:42]
  assign FPComplexAdder_io_in_a_Im = io_in_0_Im; // @[FPComplex.scala 604:42]
  assign FPComplexAdder_io_in_b_Re = io_in_1_Re; // @[FPComplex.scala 605:42]
  assign FPComplexAdder_io_in_b_Im = io_in_1_Im; // @[FPComplex.scala 605:42]
endmodule
module DFT_r_V1_nonregout(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im
);
  wire [31:0] cmplx_adj_io_in_Re; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_in_Im; // @[FFTDesigns.scala 1808:22]
  wire [7:0] cmplx_adj_io_in_adj; // @[FFTDesigns.scala 1808:22]
  wire  cmplx_adj_io_is_neg; // @[FFTDesigns.scala 1808:22]
  wire  cmplx_adj_io_is_flip; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_out_Re; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_out_Im; // @[FFTDesigns.scala 1808:22]
  wire  FPComplexMultiAdder_clock; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_reset; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_0_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_0_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_1_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_1_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_1_clock; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_1_reset; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_1_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_1_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 1839:26]
  cmplx_adj cmplx_adj ( // @[FFTDesigns.scala 1808:22]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder ( // @[FFTDesigns.scala 1839:26]
    .clock(FPComplexMultiAdder_clock),
    .reset(FPComplexMultiAdder_reset),
    .io_in_0_Re(FPComplexMultiAdder_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_io_in_1_Im),
    .io_out_Re(FPComplexMultiAdder_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_io_out_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder_1 ( // @[FFTDesigns.scala 1839:26]
    .clock(FPComplexMultiAdder_1_clock),
    .reset(FPComplexMultiAdder_1_reset),
    .io_in_0_Re(FPComplexMultiAdder_1_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_1_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_1_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_1_io_in_1_Im),
    .io_out_Re(FPComplexMultiAdder_1_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_1_io_out_Im)
  );
  assign io_out_0_Re = FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 1911:17]
  assign io_out_0_Im = FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 1911:17]
  assign io_out_1_Re = FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 1911:17]
  assign io_out_1_Im = FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 1911:17]
  assign cmplx_adj_io_in_Re = io_in_1_Re; // @[FFTDesigns.scala 1820:27]
  assign cmplx_adj_io_in_Im = io_in_1_Im; // @[FFTDesigns.scala 1820:27]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FFTDesigns.scala 1821:31]
  assign cmplx_adj_io_is_neg = 1'h1; // @[FFTDesigns.scala 1822:31]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FFTDesigns.scala 1823:32]
  assign FPComplexMultiAdder_clock = clock;
  assign FPComplexMultiAdder_reset = reset;
  assign FPComplexMultiAdder_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_1_clock = clock;
  assign FPComplexMultiAdder_1_reset = reset;
  assign FPComplexMultiAdder_1_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 1896:32]
  assign FPComplexMultiAdder_1_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 1896:32]
  assign FPComplexMultiAdder_1_io_in_1_Re = cmplx_adj_io_out_Re; // @[FFTDesigns.scala 1818:24 1824:42]
  assign FPComplexMultiAdder_1_io_in_1_Im = cmplx_adj_io_out_Im; // @[FFTDesigns.scala 1818:24 1824:42]
endmodule
module DFT_r_v2(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im
);
  wire  DFT_r_V1_nonregout_clock; // @[FFTDesigns.scala 169:24]
  wire  DFT_r_V1_nonregout_reset; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_0_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_0_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_1_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_1_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_0_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_0_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_1_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_1_Im; // @[FFTDesigns.scala 169:24]
  DFT_r_V1_nonregout DFT_r_V1_nonregout ( // @[FFTDesigns.scala 169:24]
    .clock(DFT_r_V1_nonregout_clock),
    .reset(DFT_r_V1_nonregout_reset),
    .io_in_0_Re(DFT_r_V1_nonregout_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_nonregout_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_nonregout_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_nonregout_io_in_1_Im),
    .io_out_0_Re(DFT_r_V1_nonregout_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_nonregout_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_nonregout_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_nonregout_io_out_1_Im)
  );
  assign io_out_0_Re = DFT_r_V1_nonregout_io_out_0_Re; // @[FFTDesigns.scala 171:14]
  assign io_out_0_Im = DFT_r_V1_nonregout_io_out_0_Im; // @[FFTDesigns.scala 171:14]
  assign io_out_1_Re = DFT_r_V1_nonregout_io_out_1_Re; // @[FFTDesigns.scala 171:14]
  assign io_out_1_Im = DFT_r_V1_nonregout_io_out_1_Im; // @[FFTDesigns.scala 171:14]
  assign DFT_r_V1_nonregout_clock = clock;
  assign DFT_r_V1_nonregout_reset = reset;
  assign DFT_r_V1_nonregout_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 170:15]
endmodule
module RAM_Block(
  input         clock,
  input  [2:0]  io_in_raddr,
  input  [2:0]  io_in_waddr,
  input  [31:0] io_in_data_Re,
  input  [31:0] io_in_data_Im,
  input         io_re,
  input         io_wr,
  input         io_en,
  output [31:0] io_out_data_Re,
  output [31:0] io_out_data_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_0_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Im; // @[FFTDesigns.scala 3286:18]
  wire [31:0] _GEN_33 = 3'h1 == io_in_raddr ? mem_1_Im : mem_0_Im; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_34 = 3'h2 == io_in_raddr ? mem_2_Im : _GEN_33; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_35 = 3'h3 == io_in_raddr ? mem_3_Im : _GEN_34; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_36 = 3'h4 == io_in_raddr ? mem_4_Im : _GEN_35; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_37 = 3'h5 == io_in_raddr ? mem_5_Im : _GEN_36; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_38 = 3'h6 == io_in_raddr ? mem_6_Im : _GEN_37; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_39 = 3'h7 == io_in_raddr ? mem_7_Im : _GEN_38; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_41 = 3'h1 == io_in_raddr ? mem_1_Re : mem_0_Re; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_42 = 3'h2 == io_in_raddr ? mem_2_Re : _GEN_41; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_43 = 3'h3 == io_in_raddr ? mem_3_Re : _GEN_42; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_44 = 3'h4 == io_in_raddr ? mem_4_Re : _GEN_43; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_45 = 3'h5 == io_in_raddr ? mem_5_Re : _GEN_44; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_46 = 3'h6 == io_in_raddr ? mem_6_Re : _GEN_45; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_47 = 3'h7 == io_in_raddr ? mem_7_Re : _GEN_46; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_48 = io_re ? _GEN_39 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3295:24]
  wire [31:0] _GEN_49 = io_re ? _GEN_47 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3294:24]
  assign io_out_data_Re = io_en ? _GEN_49 : 32'h0; // @[FFTDesigns.scala 3287:16 3298:22]
  assign io_out_data_Im = io_en ? _GEN_48 : 32'h0; // @[FFTDesigns.scala 3287:16 3299:22]
  always @(posedge clock) begin
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_3_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_4_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_4_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_5_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_5_Im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_6_Re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_6_Im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_7_Re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_7_Im = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PermutationModuleStreamed(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [2:0]  io_in_config_0,
  input  [2:0]  io_in_config_1,
  input  [2:0]  io_in_config_2,
  input  [2:0]  io_in_config_3,
  input  [2:0]  io_in_config_4,
  input  [2:0]  io_in_config_5,
  input  [2:0]  io_in_config_6,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
  wire  _T = io_in_config_0 == 3'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_1 = io_in_config_1 == 3'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_2 = io_in_config_2 == 3'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_3 = io_in_config_3 == 3'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_4 = io_in_config_4 == 3'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_5 = io_in_config_5 == 3'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_6 = io_in_config_6 == 3'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_8 = io_in_config_0 == 3'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_9 = io_in_config_1 == 3'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_10 = io_in_config_2 == 3'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_11 = io_in_config_3 == 3'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_12 = io_in_config_4 == 3'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_13 = io_in_config_5 == 3'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_14 = io_in_config_6 == 3'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_16 = io_in_config_0 == 3'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_17 = io_in_config_1 == 3'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_18 = io_in_config_2 == 3'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_19 = io_in_config_3 == 3'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_20 = io_in_config_4 == 3'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_21 = io_in_config_5 == 3'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_22 = io_in_config_6 == 3'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_24 = io_in_config_0 == 3'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_25 = io_in_config_1 == 3'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_26 = io_in_config_2 == 3'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_27 = io_in_config_3 == 3'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_28 = io_in_config_4 == 3'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_29 = io_in_config_5 == 3'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_30 = io_in_config_6 == 3'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_32 = io_in_config_0 == 3'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_33 = io_in_config_1 == 3'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_34 = io_in_config_2 == 3'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_35 = io_in_config_3 == 3'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_36 = io_in_config_4 == 3'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_37 = io_in_config_5 == 3'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_38 = io_in_config_6 == 3'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_40 = io_in_config_0 == 3'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_41 = io_in_config_1 == 3'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_42 = io_in_config_2 == 3'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_43 = io_in_config_3 == 3'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_44 = io_in_config_4 == 3'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_45 = io_in_config_5 == 3'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_46 = io_in_config_6 == 3'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_48 = io_in_config_0 == 3'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_49 = io_in_config_1 == 3'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_50 = io_in_config_2 == 3'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_51 = io_in_config_3 == 3'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_52 = io_in_config_4 == 3'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_53 = io_in_config_5 == 3'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_54 = io_in_config_6 == 3'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_56 = io_in_config_0 == 3'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_57 = io_in_config_1 == 3'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_58 = io_in_config_2 == 3'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_59 = io_in_config_3 == 3'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_60 = io_in_config_4 == 3'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_61 = io_in_config_5 == 3'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_62 = io_in_config_6 == 3'h7; // @[FFTDesigns.scala 3194:35]
  wire [2:0] _pms_pmx_T = _T_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_1 = _T_5 ? 3'h5 : _pms_pmx_T; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_2 = _T_4 ? 3'h4 : _pms_pmx_T_1; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_3 = _T_3 ? 3'h3 : _pms_pmx_T_2; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_4 = _T_2 ? 3'h2 : _pms_pmx_T_3; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_5 = _T_1 ? 3'h1 : _pms_pmx_T_4; // @[Mux.scala 47:70]
  wire [2:0] pms_0 = _T ? 3'h0 : _pms_pmx_T_5; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_6 = _T_14 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_7 = _T_13 ? 3'h5 : _pms_pmx_T_6; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_8 = _T_12 ? 3'h4 : _pms_pmx_T_7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_9 = _T_11 ? 3'h3 : _pms_pmx_T_8; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_10 = _T_10 ? 3'h2 : _pms_pmx_T_9; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_11 = _T_9 ? 3'h1 : _pms_pmx_T_10; // @[Mux.scala 47:70]
  wire [2:0] pms_1 = _T_8 ? 3'h0 : _pms_pmx_T_11; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_12 = _T_22 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_13 = _T_21 ? 3'h5 : _pms_pmx_T_12; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_14 = _T_20 ? 3'h4 : _pms_pmx_T_13; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_15 = _T_19 ? 3'h3 : _pms_pmx_T_14; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_16 = _T_18 ? 3'h2 : _pms_pmx_T_15; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_17 = _T_17 ? 3'h1 : _pms_pmx_T_16; // @[Mux.scala 47:70]
  wire [2:0] pms_2 = _T_16 ? 3'h0 : _pms_pmx_T_17; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_18 = _T_30 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_19 = _T_29 ? 3'h5 : _pms_pmx_T_18; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_20 = _T_28 ? 3'h4 : _pms_pmx_T_19; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_21 = _T_27 ? 3'h3 : _pms_pmx_T_20; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_22 = _T_26 ? 3'h2 : _pms_pmx_T_21; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_23 = _T_25 ? 3'h1 : _pms_pmx_T_22; // @[Mux.scala 47:70]
  wire [2:0] pms_3 = _T_24 ? 3'h0 : _pms_pmx_T_23; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_24 = _T_38 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_25 = _T_37 ? 3'h5 : _pms_pmx_T_24; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_26 = _T_36 ? 3'h4 : _pms_pmx_T_25; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_27 = _T_35 ? 3'h3 : _pms_pmx_T_26; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_28 = _T_34 ? 3'h2 : _pms_pmx_T_27; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_29 = _T_33 ? 3'h1 : _pms_pmx_T_28; // @[Mux.scala 47:70]
  wire [2:0] pms_4 = _T_32 ? 3'h0 : _pms_pmx_T_29; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_30 = _T_46 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_31 = _T_45 ? 3'h5 : _pms_pmx_T_30; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_32 = _T_44 ? 3'h4 : _pms_pmx_T_31; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_33 = _T_43 ? 3'h3 : _pms_pmx_T_32; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_34 = _T_42 ? 3'h2 : _pms_pmx_T_33; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_35 = _T_41 ? 3'h1 : _pms_pmx_T_34; // @[Mux.scala 47:70]
  wire [2:0] pms_5 = _T_40 ? 3'h0 : _pms_pmx_T_35; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_36 = _T_54 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_37 = _T_53 ? 3'h5 : _pms_pmx_T_36; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_38 = _T_52 ? 3'h4 : _pms_pmx_T_37; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_39 = _T_51 ? 3'h3 : _pms_pmx_T_38; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_40 = _T_50 ? 3'h2 : _pms_pmx_T_39; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_41 = _T_49 ? 3'h1 : _pms_pmx_T_40; // @[Mux.scala 47:70]
  wire [2:0] pms_6 = _T_48 ? 3'h0 : _pms_pmx_T_41; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_42 = _T_62 ? 3'h6 : 3'h7; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_43 = _T_61 ? 3'h5 : _pms_pmx_T_42; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_44 = _T_60 ? 3'h4 : _pms_pmx_T_43; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_45 = _T_59 ? 3'h3 : _pms_pmx_T_44; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_46 = _T_58 ? 3'h2 : _pms_pmx_T_45; // @[Mux.scala 47:70]
  wire [2:0] _pms_pmx_T_47 = _T_57 ? 3'h1 : _pms_pmx_T_46; // @[Mux.scala 47:70]
  wire [2:0] pms_7 = _T_56 ? 3'h0 : _pms_pmx_T_47; // @[Mux.scala 47:70]
  wire [31:0] _GEN_1 = 3'h1 == pms_0 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_2 = 3'h2 == pms_0 ? io_in_2_Im : _GEN_1; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_3 = 3'h3 == pms_0 ? io_in_3_Im : _GEN_2; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_4 = 3'h4 == pms_0 ? io_in_4_Im : _GEN_3; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_5 = 3'h5 == pms_0 ? io_in_5_Im : _GEN_4; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_6 = 3'h6 == pms_0 ? io_in_6_Im : _GEN_5; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_9 = 3'h1 == pms_0 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_10 = 3'h2 == pms_0 ? io_in_2_Re : _GEN_9; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_11 = 3'h3 == pms_0 ? io_in_3_Re : _GEN_10; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_12 = 3'h4 == pms_0 ? io_in_4_Re : _GEN_11; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_13 = 3'h5 == pms_0 ? io_in_5_Re : _GEN_12; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_14 = 3'h6 == pms_0 ? io_in_6_Re : _GEN_13; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_17 = 3'h1 == pms_1 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_18 = 3'h2 == pms_1 ? io_in_2_Im : _GEN_17; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_19 = 3'h3 == pms_1 ? io_in_3_Im : _GEN_18; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_20 = 3'h4 == pms_1 ? io_in_4_Im : _GEN_19; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_21 = 3'h5 == pms_1 ? io_in_5_Im : _GEN_20; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_22 = 3'h6 == pms_1 ? io_in_6_Im : _GEN_21; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_25 = 3'h1 == pms_1 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_26 = 3'h2 == pms_1 ? io_in_2_Re : _GEN_25; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_27 = 3'h3 == pms_1 ? io_in_3_Re : _GEN_26; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_28 = 3'h4 == pms_1 ? io_in_4_Re : _GEN_27; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_29 = 3'h5 == pms_1 ? io_in_5_Re : _GEN_28; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_30 = 3'h6 == pms_1 ? io_in_6_Re : _GEN_29; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_33 = 3'h1 == pms_2 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_34 = 3'h2 == pms_2 ? io_in_2_Im : _GEN_33; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_35 = 3'h3 == pms_2 ? io_in_3_Im : _GEN_34; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_36 = 3'h4 == pms_2 ? io_in_4_Im : _GEN_35; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_37 = 3'h5 == pms_2 ? io_in_5_Im : _GEN_36; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_38 = 3'h6 == pms_2 ? io_in_6_Im : _GEN_37; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_41 = 3'h1 == pms_2 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_42 = 3'h2 == pms_2 ? io_in_2_Re : _GEN_41; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_43 = 3'h3 == pms_2 ? io_in_3_Re : _GEN_42; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_44 = 3'h4 == pms_2 ? io_in_4_Re : _GEN_43; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_45 = 3'h5 == pms_2 ? io_in_5_Re : _GEN_44; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_46 = 3'h6 == pms_2 ? io_in_6_Re : _GEN_45; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_49 = 3'h1 == pms_3 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_50 = 3'h2 == pms_3 ? io_in_2_Im : _GEN_49; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_51 = 3'h3 == pms_3 ? io_in_3_Im : _GEN_50; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_52 = 3'h4 == pms_3 ? io_in_4_Im : _GEN_51; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_53 = 3'h5 == pms_3 ? io_in_5_Im : _GEN_52; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_54 = 3'h6 == pms_3 ? io_in_6_Im : _GEN_53; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_57 = 3'h1 == pms_3 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_58 = 3'h2 == pms_3 ? io_in_2_Re : _GEN_57; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_59 = 3'h3 == pms_3 ? io_in_3_Re : _GEN_58; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_60 = 3'h4 == pms_3 ? io_in_4_Re : _GEN_59; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_61 = 3'h5 == pms_3 ? io_in_5_Re : _GEN_60; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_62 = 3'h6 == pms_3 ? io_in_6_Re : _GEN_61; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_65 = 3'h1 == pms_4 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_66 = 3'h2 == pms_4 ? io_in_2_Im : _GEN_65; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_67 = 3'h3 == pms_4 ? io_in_3_Im : _GEN_66; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_68 = 3'h4 == pms_4 ? io_in_4_Im : _GEN_67; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_69 = 3'h5 == pms_4 ? io_in_5_Im : _GEN_68; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_70 = 3'h6 == pms_4 ? io_in_6_Im : _GEN_69; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_73 = 3'h1 == pms_4 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_74 = 3'h2 == pms_4 ? io_in_2_Re : _GEN_73; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_75 = 3'h3 == pms_4 ? io_in_3_Re : _GEN_74; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_76 = 3'h4 == pms_4 ? io_in_4_Re : _GEN_75; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_77 = 3'h5 == pms_4 ? io_in_5_Re : _GEN_76; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_78 = 3'h6 == pms_4 ? io_in_6_Re : _GEN_77; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_81 = 3'h1 == pms_5 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_82 = 3'h2 == pms_5 ? io_in_2_Im : _GEN_81; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_83 = 3'h3 == pms_5 ? io_in_3_Im : _GEN_82; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_84 = 3'h4 == pms_5 ? io_in_4_Im : _GEN_83; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_85 = 3'h5 == pms_5 ? io_in_5_Im : _GEN_84; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_86 = 3'h6 == pms_5 ? io_in_6_Im : _GEN_85; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_89 = 3'h1 == pms_5 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_90 = 3'h2 == pms_5 ? io_in_2_Re : _GEN_89; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_91 = 3'h3 == pms_5 ? io_in_3_Re : _GEN_90; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_92 = 3'h4 == pms_5 ? io_in_4_Re : _GEN_91; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_93 = 3'h5 == pms_5 ? io_in_5_Re : _GEN_92; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_94 = 3'h6 == pms_5 ? io_in_6_Re : _GEN_93; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_97 = 3'h1 == pms_6 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_98 = 3'h2 == pms_6 ? io_in_2_Im : _GEN_97; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_99 = 3'h3 == pms_6 ? io_in_3_Im : _GEN_98; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_100 = 3'h4 == pms_6 ? io_in_4_Im : _GEN_99; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_101 = 3'h5 == pms_6 ? io_in_5_Im : _GEN_100; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_102 = 3'h6 == pms_6 ? io_in_6_Im : _GEN_101; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_105 = 3'h1 == pms_6 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_106 = 3'h2 == pms_6 ? io_in_2_Re : _GEN_105; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_107 = 3'h3 == pms_6 ? io_in_3_Re : _GEN_106; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_108 = 3'h4 == pms_6 ? io_in_4_Re : _GEN_107; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_109 = 3'h5 == pms_6 ? io_in_5_Re : _GEN_108; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_110 = 3'h6 == pms_6 ? io_in_6_Re : _GEN_109; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_113 = 3'h1 == pms_7 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_114 = 3'h2 == pms_7 ? io_in_2_Im : _GEN_113; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_115 = 3'h3 == pms_7 ? io_in_3_Im : _GEN_114; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_116 = 3'h4 == pms_7 ? io_in_4_Im : _GEN_115; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_117 = 3'h5 == pms_7 ? io_in_5_Im : _GEN_116; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_118 = 3'h6 == pms_7 ? io_in_6_Im : _GEN_117; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_121 = 3'h1 == pms_7 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_122 = 3'h2 == pms_7 ? io_in_2_Re : _GEN_121; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_123 = 3'h3 == pms_7 ? io_in_3_Re : _GEN_122; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_124 = 3'h4 == pms_7 ? io_in_4_Re : _GEN_123; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_125 = 3'h5 == pms_7 ? io_in_5_Re : _GEN_124; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_126 = 3'h6 == pms_7 ? io_in_6_Re : _GEN_125; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_0_Re = 3'h7 == pms_0 ? io_in_7_Re : _GEN_14; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_0_Im = 3'h7 == pms_0 ? io_in_7_Im : _GEN_6; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_1_Re = 3'h7 == pms_1 ? io_in_7_Re : _GEN_30; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_1_Im = 3'h7 == pms_1 ? io_in_7_Im : _GEN_22; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_2_Re = 3'h7 == pms_2 ? io_in_7_Re : _GEN_46; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_2_Im = 3'h7 == pms_2 ? io_in_7_Im : _GEN_38; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_3_Re = 3'h7 == pms_3 ? io_in_7_Re : _GEN_62; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_3_Im = 3'h7 == pms_3 ? io_in_7_Im : _GEN_54; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_4_Re = 3'h7 == pms_4 ? io_in_7_Re : _GEN_78; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_4_Im = 3'h7 == pms_4 ? io_in_7_Im : _GEN_70; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_5_Re = 3'h7 == pms_5 ? io_in_7_Re : _GEN_94; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_5_Im = 3'h7 == pms_5 ? io_in_7_Im : _GEN_86; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_6_Re = 3'h7 == pms_6 ? io_in_7_Re : _GEN_110; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_6_Im = 3'h7 == pms_6 ? io_in_7_Im : _GEN_102; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_7_Re = 3'h7 == pms_7 ? io_in_7_Re : _GEN_126; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_7_Im = 3'h7 == pms_7 ? io_in_7_Im : _GEN_118; // @[FFTDesigns.scala 3203:{17,17}]
endmodule
module M0_Config_ROM(
  input  [1:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6,
  output [2:0] io_out_7
);
  wire [2:0] _GEN_1 = 2'h1 == io_in_cnt ? 3'h1 : 3'h0; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_cnt ? 3'h2 : _GEN_1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_cnt ? 3'h2 : 3'h1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_cnt ? 3'h3 : _GEN_5; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_9 = 2'h1 == io_in_cnt ? 3'h3 : 3'h2; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_10 = 2'h2 == io_in_cnt ? 3'h0 : _GEN_9; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_13 = 2'h1 == io_in_cnt ? 3'h0 : 3'h3; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_14 = 2'h2 == io_in_cnt ? 3'h1 : _GEN_13; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_14; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_7 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_14; // @[FFTDesigns.scala 3227:{17,17}]
endmodule
module M1_Config_ROM(
  input  [1:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6,
  output [2:0] io_out_7
);
  wire [2:0] _GEN_1 = 2'h1 == io_in_cnt ? 3'h3 : 3'h0; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_cnt ? 3'h1 : _GEN_1; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_cnt ? 3'h2 : 3'h1; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_cnt ? 3'h0 : _GEN_5; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_9 = 2'h1 == io_in_cnt ? 3'h0 : 3'h2; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_10 = 2'h2 == io_in_cnt ? 3'h3 : _GEN_9; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_13 = 2'h1 == io_in_cnt ? 3'h1 : 3'h3; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_14 = 2'h2 == io_in_cnt ? 3'h2 : _GEN_13; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_6; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_10; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_14; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_6; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_10; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_7 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_14; // @[FFTDesigns.scala 3250:{17,17}]
endmodule
module Streaming_Permute_Config(
  input  [1:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6
);
  wire [2:0] _GEN_1 = 2'h1 == io_in_cnt ? 3'h2 : 3'h0; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_cnt ? 3'h1 : _GEN_1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_cnt ? 3'h1 : 3'h2; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_cnt ? 3'h3 : _GEN_5; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_9 = 2'h1 == io_in_cnt ? 3'h3 : 3'h1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_10 = 2'h2 == io_in_cnt ? 3'h0 : _GEN_9; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_13 = 2'h1 == io_in_cnt ? 3'h0 : 3'h3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_14 = 2'h2 == io_in_cnt ? 3'h2 : _GEN_13; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_17 = 2'h1 == io_in_cnt ? 3'h6 : 3'h4; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_18 = 2'h2 == io_in_cnt ? 3'h5 : _GEN_17; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_21 = 2'h1 == io_in_cnt ? 3'h5 : 3'h6; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_22 = 2'h2 == io_in_cnt ? 3'h7 : _GEN_21; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_25 = 2'h1 == io_in_cnt ? 3'h7 : 3'h5; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_26 = 2'h2 == io_in_cnt ? 3'h4 : _GEN_25; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_6; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_10; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_14; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 3'h7 : _GEN_18; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 3'h4 : _GEN_22; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 3'h6 : _GEN_26; // @[FFTDesigns.scala 3273:{17,17}]
endmodule
module PermutationsWithStreaming(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  input         io_in_en_5,
  input         io_in_en_6,
  input         io_in_en_7,
  input         io_in_en_8,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [1:0] M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2643:27]
  wire [1:0] Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2644:29]
  reg  offset_switch; // @[FFTDesigns.scala 2627:28]
  wire [8:0] _T = {io_in_en_8,io_in_en_7,io_in_en_6,io_in_en_5,io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2628:19]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2628:26]
  reg [1:0] cnt; // @[FFTDesigns.scala 2645:22]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2649:26]
  wire [1:0] _cnt_T_1 = cnt + 2'h1; // @[FFTDesigns.scala 2651:20]
  wire  _GEN_2 = cnt == 2'h3 ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2647:32 2649:23 2652:23]
  wire [3:0] _T_6 = 3'h4 * _offset_switch_T; // @[FFTDesigns.scala 2661:54]
  wire [3:0] _GEN_110 = {{1'd0}, M0_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_8 = _GEN_110 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_9 = 3'h4 * offset_switch; // @[FFTDesigns.scala 2662:41]
  wire [3:0] _GEN_111 = {{2'd0}, cnt}; // @[FFTDesigns.scala 2662:31]
  wire [3:0] _T_11 = _GEN_111 + _T_9; // @[FFTDesigns.scala 2662:31]
  wire [3:0] _T_15 = _GEN_111 + _T_6; // @[FFTDesigns.scala 2664:31]
  wire [3:0] _GEN_113 = {{1'd0}, M1_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_18 = _GEN_113 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_114 = {{1'd0}, M0_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_22 = _GEN_114 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_117 = {{1'd0}, M1_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_32 = _GEN_117 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_118 = {{1'd0}, M0_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_36 = _GEN_118 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_121 = {{1'd0}, M1_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_46 = _GEN_121 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_122 = {{1'd0}, M0_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_50 = _GEN_122 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_125 = {{1'd0}, M1_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_60 = _GEN_125 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_126 = {{1'd0}, M0_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_64 = _GEN_126 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_129 = {{1'd0}, M1_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_74 = _GEN_129 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_130 = {{1'd0}, M0_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_78 = _GEN_130 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_133 = {{1'd0}, M1_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_88 = _GEN_133 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_134 = {{1'd0}, M0_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_92 = _GEN_134 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_137 = {{1'd0}, M1_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_102 = _GEN_137 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_138 = {{1'd0}, M0_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_106 = _GEN_138 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_141 = {{1'd0}, M1_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_116 = _GEN_141 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_6 = _T_1 ? _T_8 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_7 = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  wire [3:0] _GEN_10 = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  wire [3:0] _GEN_11 = _T_1 ? _T_18 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_19 = _T_1 ? _T_22 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_24 = _T_1 ? _T_32 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_32 = _T_1 ? _T_36 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_37 = _T_1 ? _T_46 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_45 = _T_1 ? _T_50 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_50 = _T_1 ? _T_60 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_58 = _T_1 ? _T_64 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_63 = _T_1 ? _T_74 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_71 = _T_1 ? _T_78 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_76 = _T_1 ? _T_88 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_84 = _T_1 ? _T_92 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_89 = _T_1 ? _T_102 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_97 = _T_1 ? _T_106 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_102 = _T_1 ? _T_116 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  RAM_Block RAM_Block ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block RAM_Block_1 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block RAM_Block_2 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block RAM_Block_3 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block RAM_Block_4 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block RAM_Block_5 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block RAM_Block_6 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block RAM_Block_7 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block RAM_Block_8 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block RAM_Block_9 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block RAM_Block_10 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block RAM_Block_11 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block RAM_Block_12 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block RAM_Block_13 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block RAM_Block_14 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block RAM_Block_15 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  PermutationModuleStreamed PermutationModuleStreamed ( // @[FFTDesigns.scala 2641:26]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im)
  );
  M0_Config_ROM M0_Config_ROM ( // @[FFTDesigns.scala 2642:27]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7)
  );
  M1_Config_ROM M1_Config_ROM ( // @[FFTDesigns.scala 2643:27]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7)
  );
  Streaming_Permute_Config Streaming_Permute_Config ( // @[FFTDesigns.scala 2644:29]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6)
  );
  assign io_out_0_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_0_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = _GEN_6[2:0];
  assign RAM_Block_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_io_in_data_Re = io_in_0_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_in_data_Im = io_in_0_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = _GEN_19[2:0];
  assign RAM_Block_1_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_1_io_in_data_Re = io_in_1_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_in_data_Im = io_in_1_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = _GEN_32[2:0];
  assign RAM_Block_2_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_2_io_in_data_Re = io_in_2_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_in_data_Im = io_in_2_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = _GEN_45[2:0];
  assign RAM_Block_3_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_3_io_in_data_Re = io_in_3_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_in_data_Im = io_in_3_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = _GEN_58[2:0];
  assign RAM_Block_4_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_4_io_in_data_Re = io_in_4_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_in_data_Im = io_in_4_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = _GEN_71[2:0];
  assign RAM_Block_5_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_5_io_in_data_Re = io_in_5_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_in_data_Im = io_in_5_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = _GEN_84[2:0];
  assign RAM_Block_6_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_6_io_in_data_Re = io_in_6_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_in_data_Im = io_in_6_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = _GEN_97[2:0];
  assign RAM_Block_7_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_7_io_in_data_Re = io_in_7_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_in_data_Im = io_in_7_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_8_io_in_waddr = _GEN_11[2:0];
  assign RAM_Block_8_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_8_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_9_io_in_waddr = _GEN_24[2:0];
  assign RAM_Block_9_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_9_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_10_io_in_waddr = _GEN_37[2:0];
  assign RAM_Block_10_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_10_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_11_io_in_waddr = _GEN_50[2:0];
  assign RAM_Block_11_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_11_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_12_io_in_waddr = _GEN_63[2:0];
  assign RAM_Block_12_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_12_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_13_io_in_waddr = _GEN_76[2:0];
  assign RAM_Block_13_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_13_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_14_io_in_waddr = _GEN_89[2:0];
  assign RAM_Block_14_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_14_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_15_io_in_waddr = _GEN_102[2:0];
  assign RAM_Block_15_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_15_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign M0_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2694:22]
  assign M1_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2695:22]
  assign Streaming_Permute_Config_io_in_cnt = cnt; // @[FFTDesigns.scala 2696:24]
  always @(posedge clock) begin
    offset_switch <= _T_1 & _GEN_2; // @[FFTDesigns.scala 2646:30 2691:21]
    if (reset) begin // @[FFTDesigns.scala 2645:22]
      cnt <= 2'h0; // @[FFTDesigns.scala 2645:22]
    end else if (_T_1) begin // @[FFTDesigns.scala 2646:30]
      if (cnt == 2'h3) begin // @[FFTDesigns.scala 2647:32]
        cnt <= 2'h0; // @[FFTDesigns.scala 2648:13]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2651:13]
      end
    end else begin
      cnt <= 2'h0; // @[FFTDesigns.scala 2692:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module M0_Config_ROM_1(
  input  [1:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6,
  output [2:0] io_out_7
);
  wire [2:0] _GEN_1 = 2'h1 == io_in_cnt ? 3'h1 : 3'h0; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_cnt ? 3'h2 : _GEN_1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_cnt ? 3'h2 : 3'h1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_cnt ? 3'h3 : _GEN_5; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_7 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
endmodule
module M1_Config_ROM_1(
  input  [1:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6,
  output [2:0] io_out_7
);
  wire [2:0] _GEN_1 = 2'h1 == io_in_cnt ? 3'h3 : 3'h0; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_cnt ? 3'h1 : _GEN_1; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_17 = 2'h1 == io_in_cnt ? 3'h0 : 3'h2; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_18 = 2'h2 == io_in_cnt ? 3'h3 : _GEN_17; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_18; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_18; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_18; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_7 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_18; // @[FFTDesigns.scala 3250:{17,17}]
endmodule
module Streaming_Permute_Config_1(
  input  [1:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6
);
  wire [2:0] _GEN_1 = 2'h1 == io_in_cnt ? 3'h4 : 3'h0; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_cnt ? 3'h0 : _GEN_1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_5 = 2'h1 == io_in_cnt ? 3'h0 : 3'h4; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_6 = 2'h2 == io_in_cnt ? 3'h4 : _GEN_5; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_9 = 2'h1 == io_in_cnt ? 3'h5 : 3'h1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_10 = 2'h2 == io_in_cnt ? 3'h1 : _GEN_9; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_13 = 2'h1 == io_in_cnt ? 3'h1 : 3'h5; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_14 = 2'h2 == io_in_cnt ? 3'h5 : _GEN_13; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_17 = 2'h1 == io_in_cnt ? 3'h6 : 3'h2; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_18 = 2'h2 == io_in_cnt ? 3'h2 : _GEN_17; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_21 = 2'h1 == io_in_cnt ? 3'h2 : 3'h6; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_22 = 2'h2 == io_in_cnt ? 3'h6 : _GEN_21; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_25 = 2'h1 == io_in_cnt ? 3'h7 : 3'h3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_26 = 2'h2 == io_in_cnt ? 3'h3 : _GEN_25; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 3'h4 : _GEN_2; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_6; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 3'h5 : _GEN_10; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_14; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 3'h6 : _GEN_18; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 3'h2 : _GEN_22; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 3'h7 : _GEN_26; // @[FFTDesigns.scala 3273:{17,17}]
endmodule
module PermutationsWithStreaming_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  input         io_in_en_5,
  input         io_in_en_6,
  input         io_in_en_7,
  input         io_in_en_8,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [2:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [2:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [1:0] M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2643:27]
  wire [2:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2643:27]
  wire [1:0] Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2644:29]
  reg  offset_switch; // @[FFTDesigns.scala 2627:28]
  wire [8:0] _T = {io_in_en_8,io_in_en_7,io_in_en_6,io_in_en_5,io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2628:19]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2628:26]
  reg [1:0] cnt; // @[FFTDesigns.scala 2645:22]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2649:26]
  wire [1:0] _cnt_T_1 = cnt + 2'h1; // @[FFTDesigns.scala 2651:20]
  wire  _GEN_2 = cnt == 2'h3 ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2647:32 2649:23 2652:23]
  wire [3:0] _T_6 = 3'h4 * _offset_switch_T; // @[FFTDesigns.scala 2661:54]
  wire [3:0] _GEN_110 = {{1'd0}, M0_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_8 = _GEN_110 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_9 = 3'h4 * offset_switch; // @[FFTDesigns.scala 2662:41]
  wire [3:0] _GEN_111 = {{2'd0}, cnt}; // @[FFTDesigns.scala 2662:31]
  wire [3:0] _T_11 = _GEN_111 + _T_9; // @[FFTDesigns.scala 2662:31]
  wire [3:0] _T_15 = _GEN_111 + _T_6; // @[FFTDesigns.scala 2664:31]
  wire [3:0] _GEN_113 = {{1'd0}, M1_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_18 = _GEN_113 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_114 = {{1'd0}, M0_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_22 = _GEN_114 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_117 = {{1'd0}, M1_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_32 = _GEN_117 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_118 = {{1'd0}, M0_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_36 = _GEN_118 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_121 = {{1'd0}, M1_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_46 = _GEN_121 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_122 = {{1'd0}, M0_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_50 = _GEN_122 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_125 = {{1'd0}, M1_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_60 = _GEN_125 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_126 = {{1'd0}, M0_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_64 = _GEN_126 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_129 = {{1'd0}, M1_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_74 = _GEN_129 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_130 = {{1'd0}, M0_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_78 = _GEN_130 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_133 = {{1'd0}, M1_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_88 = _GEN_133 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_134 = {{1'd0}, M0_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_92 = _GEN_134 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_137 = {{1'd0}, M1_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_102 = _GEN_137 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_138 = {{1'd0}, M0_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_106 = _GEN_138 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _GEN_141 = {{1'd0}, M1_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_116 = _GEN_141 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _GEN_6 = _T_1 ? _T_8 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_7 = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  wire [3:0] _GEN_10 = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  wire [3:0] _GEN_11 = _T_1 ? _T_18 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_19 = _T_1 ? _T_22 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_24 = _T_1 ? _T_32 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_32 = _T_1 ? _T_36 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_37 = _T_1 ? _T_46 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_45 = _T_1 ? _T_50 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_50 = _T_1 ? _T_60 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_58 = _T_1 ? _T_64 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_63 = _T_1 ? _T_74 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_71 = _T_1 ? _T_78 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_76 = _T_1 ? _T_88 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_84 = _T_1 ? _T_92 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_89 = _T_1 ? _T_102 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [3:0] _GEN_97 = _T_1 ? _T_106 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [3:0] _GEN_102 = _T_1 ? _T_116 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  RAM_Block RAM_Block ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block RAM_Block_1 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block RAM_Block_2 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block RAM_Block_3 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block RAM_Block_4 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block RAM_Block_5 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block RAM_Block_6 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block RAM_Block_7 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block RAM_Block_8 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block RAM_Block_9 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block RAM_Block_10 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block RAM_Block_11 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block RAM_Block_12 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block RAM_Block_13 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block RAM_Block_14 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block RAM_Block_15 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  PermutationModuleStreamed PermutationModuleStreamed ( // @[FFTDesigns.scala 2641:26]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im)
  );
  M0_Config_ROM_1 M0_Config_ROM ( // @[FFTDesigns.scala 2642:27]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7)
  );
  M1_Config_ROM_1 M1_Config_ROM ( // @[FFTDesigns.scala 2643:27]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7)
  );
  Streaming_Permute_Config_1 Streaming_Permute_Config ( // @[FFTDesigns.scala 2644:29]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6)
  );
  assign io_out_0_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_0_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = _GEN_6[2:0];
  assign RAM_Block_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_io_in_data_Re = io_in_0_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_in_data_Im = io_in_0_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = _GEN_19[2:0];
  assign RAM_Block_1_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_1_io_in_data_Re = io_in_1_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_in_data_Im = io_in_1_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = _GEN_32[2:0];
  assign RAM_Block_2_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_2_io_in_data_Re = io_in_2_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_in_data_Im = io_in_2_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = _GEN_45[2:0];
  assign RAM_Block_3_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_3_io_in_data_Re = io_in_3_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_in_data_Im = io_in_3_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = _GEN_58[2:0];
  assign RAM_Block_4_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_4_io_in_data_Re = io_in_4_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_in_data_Im = io_in_4_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = _GEN_71[2:0];
  assign RAM_Block_5_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_5_io_in_data_Re = io_in_5_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_in_data_Im = io_in_5_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = _GEN_84[2:0];
  assign RAM_Block_6_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_6_io_in_data_Re = io_in_6_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_in_data_Im = io_in_6_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = _GEN_97[2:0];
  assign RAM_Block_7_io_in_waddr = _GEN_7[2:0];
  assign RAM_Block_7_io_in_data_Re = io_in_7_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_in_data_Im = io_in_7_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_8_io_in_waddr = _GEN_11[2:0];
  assign RAM_Block_8_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_8_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_9_io_in_waddr = _GEN_24[2:0];
  assign RAM_Block_9_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_9_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_10_io_in_waddr = _GEN_37[2:0];
  assign RAM_Block_10_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_10_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_11_io_in_waddr = _GEN_50[2:0];
  assign RAM_Block_11_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_11_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_12_io_in_waddr = _GEN_63[2:0];
  assign RAM_Block_12_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_12_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_13_io_in_waddr = _GEN_76[2:0];
  assign RAM_Block_13_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_13_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_14_io_in_waddr = _GEN_89[2:0];
  assign RAM_Block_14_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_14_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = _GEN_10[2:0];
  assign RAM_Block_15_io_in_waddr = _GEN_102[2:0];
  assign RAM_Block_15_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_15_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign M0_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2694:22]
  assign M1_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2695:22]
  assign Streaming_Permute_Config_io_in_cnt = cnt; // @[FFTDesigns.scala 2696:24]
  always @(posedge clock) begin
    offset_switch <= _T_1 & _GEN_2; // @[FFTDesigns.scala 2646:30 2691:21]
    if (reset) begin // @[FFTDesigns.scala 2645:22]
      cnt <= 2'h0; // @[FFTDesigns.scala 2645:22]
    end else if (_T_1) begin // @[FFTDesigns.scala 2646:30]
      if (cnt == 2'h3) begin // @[FFTDesigns.scala 2647:32]
        cnt <= 2'h0; // @[FFTDesigns.scala 2648:13]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2651:13]
      end
    end else begin
      cnt <= 2'h0; // @[FFTDesigns.scala 2692:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM(
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im
);
  wire [31:0] _GEN_10 = 2'h2 == io_in_addr[1:0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_14 = 2'h2 == io_in_addr[1:0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_1_Re = 2'h3 == io_in_addr[1:0] ? 32'h248d3131 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_1_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_3_Re = 2'h3 == io_in_addr[1:0] ? 32'h248d3131 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_3_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_5_Re = 2'h3 == io_in_addr[1:0] ? 32'h248d3131 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_5_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_7_Re = 2'h3 == io_in_addr[1:0] ? 32'h248d3131 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_7_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
endmodule
module TwiddleFactorsStreamed(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] TwiddleFactorROM_io_in_addr; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] cmplx_adj_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_1_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_1_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_1_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_1_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_1_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_1_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_1_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_2_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_2_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_2_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_2_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_2_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_2_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_2_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_3_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_3_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_3_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_3_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_3_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_3_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_3_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_4_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_4_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_4_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_4_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_4_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_4_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_4_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_5_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_5_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_5_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_5_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_5_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_5_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_5_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_6_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_6_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_6_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_6_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_6_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_6_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_6_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_7_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_7_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_7_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_7_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_7_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_7_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_7_io_out_Im; // @[FFTDesigns.scala 2146:30]
  reg [1:0] cnt; // @[FFTDesigns.scala 2139:24]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2140:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2140:28]
  wire [1:0] _cnt_T_1 = cnt + 2'h1; // @[FFTDesigns.scala 2153:22]
  wire  _GEN_8 = TwiddleFactorROM_io_out_data_1_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_9 = TwiddleFactorROM_io_out_data_1_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_1_Re[31] :
    TwiddleFactorROM_io_out_data_1_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_16 = TwiddleFactorROM_io_out_data_3_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_17 = TwiddleFactorROM_io_out_data_3_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_3_Re[31] :
    TwiddleFactorROM_io_out_data_3_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_24 = TwiddleFactorROM_io_out_data_5_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_25 = TwiddleFactorROM_io_out_data_5_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_5_Re[31] :
    TwiddleFactorROM_io_out_data_5_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_32 = TwiddleFactorROM_io_out_data_7_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_33 = TwiddleFactorROM_io_out_data_7_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_7_Re[31] :
    TwiddleFactorROM_io_out_data_7_Im[31]; // @[FFTDesigns.scala 2158:92]
  reg [31:0] result_regs_0_0_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_0_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_1_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_1_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_2_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_2_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_3_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_3_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_4_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_4_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_5_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_5_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_6_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_6_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_7_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_7_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_0_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_0_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_1_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_1_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_2_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_2_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_3_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_3_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_4_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_4_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_5_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_5_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_6_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_6_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_7_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_7_Im; // @[FFTDesigns.scala 2183:32]
  TwiddleFactorROM TwiddleFactorROM ( // @[FFTDesigns.scala 2098:26]
    .io_in_addr(TwiddleFactorROM_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_io_out_data_1_Im),
    .io_out_data_3_Re(TwiddleFactorROM_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_io_out_data_3_Im),
    .io_out_data_5_Re(TwiddleFactorROM_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_io_out_data_7_Im)
  );
  cmplx_adj cmplx_adj ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  cmplx_adj cmplx_adj_1 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_1_io_in_Re),
    .io_in_Im(cmplx_adj_1_io_in_Im),
    .io_in_adj(cmplx_adj_1_io_in_adj),
    .io_is_neg(cmplx_adj_1_io_is_neg),
    .io_is_flip(cmplx_adj_1_io_is_flip),
    .io_out_Re(cmplx_adj_1_io_out_Re),
    .io_out_Im(cmplx_adj_1_io_out_Im)
  );
  cmplx_adj cmplx_adj_2 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_2_io_in_Re),
    .io_in_Im(cmplx_adj_2_io_in_Im),
    .io_in_adj(cmplx_adj_2_io_in_adj),
    .io_is_neg(cmplx_adj_2_io_is_neg),
    .io_is_flip(cmplx_adj_2_io_is_flip),
    .io_out_Re(cmplx_adj_2_io_out_Re),
    .io_out_Im(cmplx_adj_2_io_out_Im)
  );
  cmplx_adj cmplx_adj_3 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_3_io_in_Re),
    .io_in_Im(cmplx_adj_3_io_in_Im),
    .io_in_adj(cmplx_adj_3_io_in_adj),
    .io_is_neg(cmplx_adj_3_io_is_neg),
    .io_is_flip(cmplx_adj_3_io_is_flip),
    .io_out_Re(cmplx_adj_3_io_out_Re),
    .io_out_Im(cmplx_adj_3_io_out_Im)
  );
  cmplx_adj cmplx_adj_4 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_4_io_in_Re),
    .io_in_Im(cmplx_adj_4_io_in_Im),
    .io_in_adj(cmplx_adj_4_io_in_adj),
    .io_is_neg(cmplx_adj_4_io_is_neg),
    .io_is_flip(cmplx_adj_4_io_is_flip),
    .io_out_Re(cmplx_adj_4_io_out_Re),
    .io_out_Im(cmplx_adj_4_io_out_Im)
  );
  cmplx_adj cmplx_adj_5 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_5_io_in_Re),
    .io_in_Im(cmplx_adj_5_io_in_Im),
    .io_in_adj(cmplx_adj_5_io_in_adj),
    .io_is_neg(cmplx_adj_5_io_is_neg),
    .io_is_flip(cmplx_adj_5_io_is_flip),
    .io_out_Re(cmplx_adj_5_io_out_Re),
    .io_out_Im(cmplx_adj_5_io_out_Im)
  );
  cmplx_adj cmplx_adj_6 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_6_io_in_Re),
    .io_in_Im(cmplx_adj_6_io_in_Im),
    .io_in_adj(cmplx_adj_6_io_in_adj),
    .io_is_neg(cmplx_adj_6_io_is_neg),
    .io_is_flip(cmplx_adj_6_io_is_flip),
    .io_out_Re(cmplx_adj_6_io_out_Re),
    .io_out_Im(cmplx_adj_6_io_out_Im)
  );
  cmplx_adj cmplx_adj_7 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_7_io_in_Re),
    .io_in_Im(cmplx_adj_7_io_in_Im),
    .io_in_adj(cmplx_adj_7_io_in_adj),
    .io_is_neg(cmplx_adj_7_io_is_neg),
    .io_is_flip(cmplx_adj_7_io_is_flip),
    .io_out_Re(cmplx_adj_7_io_out_Re),
    .io_out_Im(cmplx_adj_7_io_out_Im)
  );
  assign io_out_0_Re = result_regs_1_0_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_0_Im = result_regs_1_0_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_1_Re = result_regs_1_1_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_1_Im = result_regs_1_1_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_2_Re = result_regs_1_2_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_2_Im = result_regs_1_2_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_3_Re = result_regs_1_3_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_3_Im = result_regs_1_3_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_4_Re = result_regs_1_4_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_4_Im = result_regs_1_4_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_5_Re = result_regs_1_5_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_5_Im = result_regs_1_5_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_6_Re = result_regs_1_6_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_6_Im = result_regs_1_6_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_7_Re = result_regs_1_7_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_7_Im = result_regs_1_7_Im; // @[FFTDesigns.scala 2193:14]
  assign TwiddleFactorROM_io_in_addr = {{3'd0}, cnt}; // @[FFTDesigns.scala 2194:24]
  assign cmplx_adj_io_in_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_io_in_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_io_in_adj = 8'h0;
  assign cmplx_adj_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_1_io_in_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_1_io_in_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_1_io_in_adj = 8'h0;
  assign cmplx_adj_1_io_is_neg = _T_1 & _GEN_9; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_1_io_is_flip = _T_1 & _GEN_8; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_2_io_in_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_2_io_in_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_2_io_in_adj = 8'h0;
  assign cmplx_adj_2_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_2_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_3_io_in_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_3_io_in_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_3_io_in_adj = 8'h0;
  assign cmplx_adj_3_io_is_neg = _T_1 & _GEN_17; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_3_io_is_flip = _T_1 & _GEN_16; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_4_io_in_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_4_io_in_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_4_io_in_adj = 8'h0;
  assign cmplx_adj_4_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_4_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_5_io_in_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_5_io_in_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_5_io_in_adj = 8'h0;
  assign cmplx_adj_5_io_is_neg = _T_1 & _GEN_25; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_5_io_is_flip = _T_1 & _GEN_24; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_6_io_in_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_6_io_in_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_6_io_in_adj = 8'h0;
  assign cmplx_adj_6_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_6_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_7_io_in_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_7_io_in_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_7_io_in_adj = 8'h0;
  assign cmplx_adj_7_io_is_neg = _T_1 & _GEN_33; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_7_io_is_flip = _T_1 & _GEN_32; // @[FFTDesigns.scala 2149:32 2179:34]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2139:24]
      cnt <= 2'h0; // @[FFTDesigns.scala 2139:24]
    end else if (_T_1) begin // @[FFTDesigns.scala 2149:32]
      if (cnt == 2'h3) begin // @[FFTDesigns.scala 2150:34]
        cnt <= 2'h0; // @[FFTDesigns.scala 2151:15]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2153:15]
      end
    end else begin
      cnt <= 2'h0; // @[FFTDesigns.scala 2175:13]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_0_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_0_Re <= cmplx_adj_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_0_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_0_Im <= cmplx_adj_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_1_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_1_Re <= cmplx_adj_1_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_1_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_1_Im <= cmplx_adj_1_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_2_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_2_Re <= cmplx_adj_2_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_2_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_2_Im <= cmplx_adj_2_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_3_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_3_Re <= cmplx_adj_3_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_3_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_3_Im <= cmplx_adj_3_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_4_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_4_Re <= cmplx_adj_4_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_4_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_4_Im <= cmplx_adj_4_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_5_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_5_Re <= cmplx_adj_5_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_5_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_5_Im <= cmplx_adj_5_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_6_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_6_Re <= cmplx_adj_6_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_6_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_6_Im <= cmplx_adj_6_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_7_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_7_Re <= cmplx_adj_7_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_7_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_7_Im <= cmplx_adj_7_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_0_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_0_Re <= result_regs_0_0_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_0_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_0_Im <= result_regs_0_0_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_1_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_1_Re <= result_regs_0_1_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_1_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_1_Im <= result_regs_0_1_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_2_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_2_Re <= result_regs_0_2_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_2_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_2_Im <= result_regs_0_2_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_3_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_3_Re <= result_regs_0_3_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_3_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_3_Im <= result_regs_0_3_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_4_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_4_Re <= result_regs_0_4_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_4_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_4_Im <= result_regs_0_4_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_5_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_5_Re <= result_regs_0_5_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_5_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_5_Im <= result_regs_0_5_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_6_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_6_Re <= result_regs_0_6_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_6_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_6_Im <= result_regs_0_6_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_7_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_7_Re <= result_regs_0_7_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_7_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_7_Im <= result_regs_0_7_Im; // @[FFTDesigns.scala 2190:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  result_regs_0_0_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  result_regs_0_0_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  result_regs_0_1_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  result_regs_0_1_Im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  result_regs_0_2_Re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  result_regs_0_2_Im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  result_regs_0_3_Re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  result_regs_0_3_Im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  result_regs_0_4_Re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  result_regs_0_4_Im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  result_regs_0_5_Re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  result_regs_0_5_Im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  result_regs_0_6_Re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  result_regs_0_6_Im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  result_regs_0_7_Re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  result_regs_0_7_Im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  result_regs_1_0_Re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  result_regs_1_0_Im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  result_regs_1_1_Re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  result_regs_1_1_Im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  result_regs_1_2_Re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  result_regs_1_2_Im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  result_regs_1_3_Re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  result_regs_1_3_Im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  result_regs_1_4_Re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  result_regs_1_4_Im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  result_regs_1_5_Re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  result_regs_1_5_Im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  result_regs_1_6_Re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  result_regs_1_6_Im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  result_regs_1_7_Re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  result_regs_1_7_Im = _RAND_32[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_1(
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im
);
  wire [31:0] _GEN_9 = 2'h1 == io_in_addr[1:0] ? 32'h3f3504f2 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_10 = 2'h2 == io_in_addr[1:0] ? 32'h248d3131 : _GEN_9; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_13 = 2'h1 == io_in_addr[1:0] ? 32'hbf3504f2 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_14 = 2'h2 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_13; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_1_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_1_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_3_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_3_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_5_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_5_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_7_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_7_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
endmodule
module FP_subber(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_clock; // @[FPArithmetic.scala 414:26]
  wire  FP_adder_reset; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_in_a; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_in_b; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_out_s; // @[FPArithmetic.scala 414:26]
  wire  _adjusted_in_b_T_1 = ~io_in_b[31]; // @[FPArithmetic.scala 417:23]
  FP_adder FP_adder ( // @[FPArithmetic.scala 414:26]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  assign io_out_s = FP_adder_io_out_s; // @[FPArithmetic.scala 420:14]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = io_in_a; // @[FPArithmetic.scala 418:22]
  assign FP_adder_io_in_b = {_adjusted_in_b_T_1,io_in_b[30:0]}; // @[FPArithmetic.scala 417:39]
endmodule
module multiplier(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[Arithmetic.scala 84:23]
endmodule
module full_adder_82(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 58:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 58:34]
  wire [8:0] result = _result_T_1[8:0]; // @[Arithmetic.scala 57:22 58:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 59:23]
endmodule
module FP_multiplier(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] multiplier_io_in_a; // @[FPArithmetic.scala 488:28]
  wire [23:0] multiplier_io_in_b; // @[FPArithmetic.scala 488:28]
  wire [47:0] multiplier_io_out_s; // @[FPArithmetic.scala 488:28]
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 493:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 493:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 493:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 493:24]
  wire [7:0] complementN_io_in; // @[FPArithmetic.scala 499:29]
  wire [7:0] complementN_io_out; // @[FPArithmetic.scala 499:29]
  wire [7:0] adderN_io_in_a; // @[FPArithmetic.scala 503:24]
  wire [7:0] adderN_io_in_b; // @[FPArithmetic.scala 503:24]
  wire [7:0] adderN_io_out_s; // @[FPArithmetic.scala 503:24]
  wire  s_0 = io_in_a[31]; // @[FPArithmetic.scala 453:20]
  wire  s_1 = io_in_b[31]; // @[FPArithmetic.scala 454:20]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 458:62]
  wire [8:0] _GEN_13 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 458:34]
  wire [8:0] _GEN_0 = _GEN_13 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 458:68 459:14 461:14]
  wire [8:0] _GEN_14 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 463:34]
  wire [8:0] _GEN_1 = _GEN_14 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 463:68 464:14 466:14]
  wire [22:0] exp_check_0 = {{15'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 469:25 470:18]
  wire [22:0] _cond_holder_T_1 = exp_check_0 + 23'h1; // @[FPArithmetic.scala 474:34]
  wire [22:0] exp_check_1 = {{15'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 469:25 471:18]
  wire [22:0] _cond_holder_T_3 = 23'h7f - exp_check_1; // @[FPArithmetic.scala 474:80]
  wire [22:0] _cond_holder_T_4 = ~_cond_holder_T_3; // @[FPArithmetic.scala 474:42]
  wire [22:0] _cond_holder_T_6 = _cond_holder_T_1 + _cond_holder_T_4; // @[FPArithmetic.scala 474:40]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 478:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 479:23]
  wire  new_s = s_0 ^ s_1; // @[FPArithmetic.scala 510:19]
  wire [7:0] _new_exp_T_1 = adderN_io_out_s + 8'h1; // @[FPArithmetic.scala 521:34]
  wire [22:0] _cond_holder_T_8 = exp_check_0 + 23'h2; // @[FPArithmetic.scala 523:36]
  wire [22:0] _cond_holder_T_13 = _cond_holder_T_8 + _cond_holder_T_4; // @[FPArithmetic.scala 523:42]
  wire [23:0] _new_mant_T_2 = {multiplier_io_out_s[46:24], 1'h0}; // @[FPArithmetic.scala 529:73]
  wire [7:0] _GEN_2 = multiplier_io_out_s[47] ? _new_exp_T_1 : adderN_io_out_s; // @[FPArithmetic.scala 520:60 521:15 526:15]
  wire [22:0] cond_holder = multiplier_io_out_s[47] ? _cond_holder_T_13 : _cond_holder_T_6; // @[FPArithmetic.scala 520:60 523:19 528:19]
  wire [23:0] _GEN_5 = multiplier_io_out_s[47] ? {{1'd0}, multiplier_io_out_s[46:24]} : _new_mant_T_2; // @[FPArithmetic.scala 520:60 524:16 529:16]
  reg [31:0] reg_out_s; // @[FPArithmetic.scala 531:28]
  wire [22:0] _T_12 = ~cond_holder; // @[FPArithmetic.scala 533:51]
  wire [22:0] _T_14 = 23'h1 + _T_12; // @[FPArithmetic.scala 533:49]
  wire [22:0] _GEN_15 = {{14'd0}, _T_2}; // @[FPArithmetic.scala 533:42]
  wire [8:0] _GEN_6 = cond_holder > _GEN_15 ? _T_2 : {{1'd0}, _GEN_2}; // @[FPArithmetic.scala 538:61 539:15]
  wire [8:0] _GEN_9 = _GEN_15 >= _T_14 ? 9'h1 : _GEN_6; // @[FPArithmetic.scala 533:67 534:15]
  wire [7:0] new_exp = _GEN_9[7:0]; // @[FPArithmetic.scala 513:23]
  wire [23:0] _new_mant_T_4 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 540:45]
  wire [23:0] _GEN_7 = cond_holder > _GEN_15 ? _new_mant_T_4 : _GEN_5; // @[FPArithmetic.scala 538:61 540:16]
  wire [23:0] _GEN_10 = _GEN_15 >= _T_14 ? 24'h400000 : _GEN_7; // @[FPArithmetic.scala 533:67 535:16]
  wire [22:0] new_mant = _GEN_10[22:0]; // @[FPArithmetic.scala 515:24]
  wire [31:0] _reg_out_s_T_1 = {new_s,new_exp,new_mant}; // @[FPArithmetic.scala 536:37]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 457:19]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 457:19]
  multiplier multiplier ( // @[FPArithmetic.scala 488:28]
    .io_in_a(multiplier_io_in_a),
    .io_in_b(multiplier_io_in_b),
    .io_out_s(multiplier_io_out_s)
  );
  full_subber subber ( // @[FPArithmetic.scala 493:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complementN ( // @[FPArithmetic.scala 499:29]
    .io_in(complementN_io_in),
    .io_out(complementN_io_out)
  );
  full_adder_82 adderN ( // @[FPArithmetic.scala 503:24]
    .io_in_a(adderN_io_in_a),
    .io_in_b(adderN_io_in_b),
    .io_out_s(adderN_io_out_s)
  );
  assign io_out_s = reg_out_s; // @[FPArithmetic.scala 548:14]
  assign multiplier_io_in_a = {1'h1,frac_0}; // @[FPArithmetic.scala 483:24]
  assign multiplier_io_in_b = {1'h1,frac_1}; // @[FPArithmetic.scala 484:24]
  assign subber_io_in_a = 8'h7f; // @[FPArithmetic.scala 494:20]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 457:19]
  assign complementN_io_in = subber_io_out_s; // @[FPArithmetic.scala 500:23]
  assign adderN_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 457:19]
  assign adderN_io_in_b = complementN_io_out; // @[FPArithmetic.scala 505:20]
  always @(posedge clock) begin
    if (reset) begin // @[FPArithmetic.scala 531:28]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 531:28]
    end else if (exp_0 == 8'h0 | exp_1 == 8'h0) begin // @[FPArithmetic.scala 543:43]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 544:17]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FPArithmetic.scala 546:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_out_s = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMult(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_subber_clock; // @[FPComplex.scala 123:24]
  wire  FP_subber_reset; // @[FPComplex.scala 123:24]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 123:24]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 123:24]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 123:24]
  wire  FP_adder_clock; // @[FPComplex.scala 124:24]
  wire  FP_adder_reset; // @[FPComplex.scala 124:24]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 124:24]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 124:24]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 124:24]
  wire  FP_multiplier_clock; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_reset; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_1_reset; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_2_clock; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_2_reset; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_2_io_in_a; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_2_io_in_b; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_2_io_out_s; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_3_clock; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_3_reset; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_3_io_in_a; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_3_io_in_b; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_3_io_out_s; // @[FPComplex.scala 126:26]
  FP_subber FP_subber ( // @[FPComplex.scala 123:24]
    .clock(FP_subber_clock),
    .reset(FP_subber_reset),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_adder FP_adder ( // @[FPComplex.scala 124:24]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 126:26]
    .clock(FP_multiplier_clock),
    .reset(FP_multiplier_reset),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 126:26]
    .clock(FP_multiplier_1_clock),
    .reset(FP_multiplier_1_reset),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  FP_multiplier FP_multiplier_2 ( // @[FPComplex.scala 126:26]
    .clock(FP_multiplier_2_clock),
    .reset(FP_multiplier_2_reset),
    .io_in_a(FP_multiplier_2_io_in_a),
    .io_in_b(FP_multiplier_2_io_in_b),
    .io_out_s(FP_multiplier_2_io_out_s)
  );
  FP_multiplier FP_multiplier_3 ( // @[FPComplex.scala 126:26]
    .clock(FP_multiplier_3_clock),
    .reset(FP_multiplier_3_reset),
    .io_in_a(FP_multiplier_3_io_in_a),
    .io_in_b(FP_multiplier_3_io_in_b),
    .io_out_s(FP_multiplier_3_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 141:17]
  assign io_out_s_Im = FP_adder_io_out_s; // @[FPComplex.scala 142:17]
  assign FP_subber_clock = clock;
  assign FP_subber_reset = reset;
  assign FP_subber_io_in_a = FP_multiplier_io_out_s; // @[FPComplex.scala 137:17]
  assign FP_subber_io_in_b = FP_multiplier_1_io_out_s; // @[FPComplex.scala 138:17]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = FP_multiplier_2_io_out_s; // @[FPComplex.scala 139:17]
  assign FP_adder_io_in_b = FP_multiplier_3_io_out_s; // @[FPComplex.scala 140:17]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_reset = reset;
  assign FP_multiplier_io_in_a = io_in_a_Re; // @[FPComplex.scala 129:28]
  assign FP_multiplier_io_in_b = io_in_b_Re; // @[FPComplex.scala 130:28]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_reset = reset;
  assign FP_multiplier_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 131:28]
  assign FP_multiplier_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 132:28]
  assign FP_multiplier_2_clock = clock;
  assign FP_multiplier_2_reset = reset;
  assign FP_multiplier_2_io_in_a = io_in_a_Re; // @[FPComplex.scala 133:28]
  assign FP_multiplier_2_io_in_b = io_in_b_Im; // @[FPComplex.scala 134:28]
  assign FP_multiplier_3_clock = clock;
  assign FP_multiplier_3_reset = reset;
  assign FP_multiplier_3_io_in_a = io_in_a_Im; // @[FPComplex.scala 135:28]
  assign FP_multiplier_3_io_in_b = io_in_b_Re; // @[FPComplex.scala 136:28]
endmodule
module TwiddleFactorsStreamed_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] TwiddleFactorROM_io_in_addr; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Im; // @[FFTDesigns.scala 2098:26]
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  reg [1:0] cnt; // @[FFTDesigns.scala 2106:24]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2107:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2107:28]
  wire [1:0] _cnt_T_1 = cnt + 2'h1; // @[FFTDesigns.scala 2120:22]
  TwiddleFactorROM_1 TwiddleFactorROM ( // @[FFTDesigns.scala 2098:26]
    .io_in_addr(TwiddleFactorROM_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_io_out_data_1_Im),
    .io_out_data_3_Re(TwiddleFactorROM_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_io_out_data_3_Im),
    .io_out_data_5_Re(TwiddleFactorROM_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_io_out_data_7_Im)
  );
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_clock),
    .reset(FPComplexMult_reset),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_1_clock),
    .reset(FPComplexMult_1_reset),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_2_clock),
    .reset(FPComplexMult_2_reset),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_3_clock),
    .reset(FPComplexMult_3_reset),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_4_clock),
    .reset(FPComplexMult_4_reset),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_5_clock),
    .reset(FPComplexMult_5_reset),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_6_clock),
    .reset(FPComplexMult_6_reset),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_7_clock),
    .reset(FPComplexMult_7_reset),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign TwiddleFactorROM_io_in_addr = {{3'd0}, cnt}; // @[FFTDesigns.scala 2136:24]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_reset = reset;
  assign FPComplexMult_io_in_a_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_a_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_reset = reset;
  assign FPComplexMult_1_io_in_a_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_a_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_reset = reset;
  assign FPComplexMult_2_io_in_a_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_a_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_reset = reset;
  assign FPComplexMult_3_io_in_a_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_a_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_reset = reset;
  assign FPComplexMult_4_io_in_a_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_a_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_reset = reset;
  assign FPComplexMult_5_io_in_a_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_a_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_reset = reset;
  assign FPComplexMult_6_io_in_a_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_a_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_reset = reset;
  assign FPComplexMult_7_io_in_a_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_a_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2106:24]
      cnt <= 2'h0; // @[FFTDesigns.scala 2106:24]
    end else if (_T_1) begin // @[FFTDesigns.scala 2116:32]
      if (cnt == 2'h3) begin // @[FFTDesigns.scala 2117:34]
        cnt <= 2'h0; // @[FFTDesigns.scala 2118:15]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2120:15]
      end
    end else begin
      cnt <= 2'h0; // @[FFTDesigns.scala 2131:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_2(
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im
);
  wire [31:0] _GEN_9 = 2'h1 == io_in_addr[1:0] ? 32'h3f3504f2 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_10 = 2'h2 == io_in_addr[1:0] ? 32'h248d3131 : _GEN_9; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_13 = 2'h1 == io_in_addr[1:0] ? 32'hbf3504f2 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_14 = 2'h2 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_13; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_41 = 2'h1 == io_in_addr[1:0] ? 32'h3ec3ef14 : 32'h3f6c835e; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_42 = 2'h2 == io_in_addr[1:0] ? 32'hbec3ef14 : _GEN_41; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_45 = 2'h1 == io_in_addr[1:0] ? 32'hbf6c835e : 32'hbec3ef14; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_46 = 2'h2 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_45; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_1_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_1_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_3_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_3_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_5_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_42; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_5_Im = 2'h3 == io_in_addr[1:0] ? 32'hbec3ef14 : _GEN_46; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_7_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_42; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_7_Im = 2'h3 == io_in_addr[1:0] ? 32'hbec3ef14 : _GEN_46; // @[FFTDesigns.scala 2059:{25,25}]
endmodule
module TwiddleFactorsStreamed_2(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] TwiddleFactorROM_io_in_addr; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Im; // @[FFTDesigns.scala 2098:26]
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  reg [1:0] cnt; // @[FFTDesigns.scala 2106:24]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2107:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2107:28]
  wire [1:0] _cnt_T_1 = cnt + 2'h1; // @[FFTDesigns.scala 2120:22]
  TwiddleFactorROM_2 TwiddleFactorROM ( // @[FFTDesigns.scala 2098:26]
    .io_in_addr(TwiddleFactorROM_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_io_out_data_1_Im),
    .io_out_data_3_Re(TwiddleFactorROM_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_io_out_data_3_Im),
    .io_out_data_5_Re(TwiddleFactorROM_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_io_out_data_7_Im)
  );
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_clock),
    .reset(FPComplexMult_reset),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_1_clock),
    .reset(FPComplexMult_1_reset),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_2_clock),
    .reset(FPComplexMult_2_reset),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_3_clock),
    .reset(FPComplexMult_3_reset),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_4_clock),
    .reset(FPComplexMult_4_reset),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_5_clock),
    .reset(FPComplexMult_5_reset),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_6_clock),
    .reset(FPComplexMult_6_reset),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_7_clock),
    .reset(FPComplexMult_7_reset),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign TwiddleFactorROM_io_in_addr = {{3'd0}, cnt}; // @[FFTDesigns.scala 2136:24]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_reset = reset;
  assign FPComplexMult_io_in_a_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_a_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_reset = reset;
  assign FPComplexMult_1_io_in_a_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_a_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_reset = reset;
  assign FPComplexMult_2_io_in_a_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_a_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_reset = reset;
  assign FPComplexMult_3_io_in_a_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_a_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_reset = reset;
  assign FPComplexMult_4_io_in_a_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_a_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_reset = reset;
  assign FPComplexMult_5_io_in_a_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_a_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_reset = reset;
  assign FPComplexMult_6_io_in_a_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_a_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_reset = reset;
  assign FPComplexMult_7_io_in_a_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_a_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2106:24]
      cnt <= 2'h0; // @[FFTDesigns.scala 2106:24]
    end else if (_T_1) begin // @[FFTDesigns.scala 2116:32]
      if (cnt == 2'h3) begin // @[FFTDesigns.scala 2117:34]
        cnt <= 2'h0; // @[FFTDesigns.scala 2118:15]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2120:15]
      end
    end else begin
      cnt <= 2'h0; // @[FFTDesigns.scala 2131:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_3(
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im
);
  wire [31:0] _GEN_9 = 2'h1 == io_in_addr[1:0] ? 32'h3f3504f2 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_10 = 2'h2 == io_in_addr[1:0] ? 32'h248d3131 : _GEN_9; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_13 = 2'h1 == io_in_addr[1:0] ? 32'hbf3504f2 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_14 = 2'h2 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_13; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_25 = 2'h1 == io_in_addr[1:0] ? 32'h3f0e39d8 : 32'h3f7b14be; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_26 = 2'h2 == io_in_addr[1:0] ? 32'hbe47c5c0 : _GEN_25; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_29 = 2'h1 == io_in_addr[1:0] ? 32'hbf54db30 : 32'hbe47c5c0; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_30 = 2'h2 == io_in_addr[1:0] ? 32'hbf7b14be : _GEN_29; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_41 = 2'h1 == io_in_addr[1:0] ? 32'h3ec3ef14 : 32'h3f6c835e; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_42 = 2'h2 == io_in_addr[1:0] ? 32'hbec3ef14 : _GEN_41; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_45 = 2'h1 == io_in_addr[1:0] ? 32'hbf6c835e : 32'hbec3ef14; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_46 = 2'h2 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_45; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_57 = 2'h1 == io_in_addr[1:0] ? 32'h3e47c5c0 : 32'h3f54db30; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_58 = 2'h2 == io_in_addr[1:0] ? 32'hbf0e39d8 : _GEN_57; // @[FFTDesigns.scala 2058:{25,25}]
  wire [31:0] _GEN_61 = 2'h1 == io_in_addr[1:0] ? 32'hbf7b14be : 32'hbf0e39d8; // @[FFTDesigns.scala 2059:{25,25}]
  wire [31:0] _GEN_62 = 2'h2 == io_in_addr[1:0] ? 32'hbf54db30 : _GEN_61; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_1_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_10; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_1_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_3_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf54db30 : _GEN_26; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_3_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf0e39d8 : _GEN_30; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_5_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_42; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_5_Im = 2'h3 == io_in_addr[1:0] ? 32'hbec3ef14 : _GEN_46; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_7_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf7b14be : _GEN_58; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_7_Im = 2'h3 == io_in_addr[1:0] ? 32'hbe47c5c0 : _GEN_62; // @[FFTDesigns.scala 2059:{25,25}]
endmodule
module TwiddleFactorsStreamed_3(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] TwiddleFactorROM_io_in_addr; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Im; // @[FFTDesigns.scala 2098:26]
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  reg [1:0] cnt; // @[FFTDesigns.scala 2106:24]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2107:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2107:28]
  wire [1:0] _cnt_T_1 = cnt + 2'h1; // @[FFTDesigns.scala 2120:22]
  TwiddleFactorROM_3 TwiddleFactorROM ( // @[FFTDesigns.scala 2098:26]
    .io_in_addr(TwiddleFactorROM_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_io_out_data_1_Im),
    .io_out_data_3_Re(TwiddleFactorROM_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_io_out_data_3_Im),
    .io_out_data_5_Re(TwiddleFactorROM_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_io_out_data_7_Im)
  );
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_clock),
    .reset(FPComplexMult_reset),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_1_clock),
    .reset(FPComplexMult_1_reset),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_2_clock),
    .reset(FPComplexMult_2_reset),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_3_clock),
    .reset(FPComplexMult_3_reset),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_4_clock),
    .reset(FPComplexMult_4_reset),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_5_clock),
    .reset(FPComplexMult_5_reset),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_6_clock),
    .reset(FPComplexMult_6_reset),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_7_clock),
    .reset(FPComplexMult_7_reset),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign TwiddleFactorROM_io_in_addr = {{3'd0}, cnt}; // @[FFTDesigns.scala 2136:24]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_reset = reset;
  assign FPComplexMult_io_in_a_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_a_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_reset = reset;
  assign FPComplexMult_1_io_in_a_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_a_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_reset = reset;
  assign FPComplexMult_2_io_in_a_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_a_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_reset = reset;
  assign FPComplexMult_3_io_in_a_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_a_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_reset = reset;
  assign FPComplexMult_4_io_in_a_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_a_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_reset = reset;
  assign FPComplexMult_5_io_in_a_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_a_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_reset = reset;
  assign FPComplexMult_6_io_in_a_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_a_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_reset = reset;
  assign FPComplexMult_7_io_in_a_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_a_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2106:24]
      cnt <= 2'h0; // @[FFTDesigns.scala 2106:24]
    end else if (_T_1) begin // @[FFTDesigns.scala 2116:32]
      if (cnt == 2'h3) begin // @[FFTDesigns.scala 2117:34]
        cnt <= 2'h0; // @[FFTDesigns.scala 2118:15]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2120:15]
      end
    end else begin
      cnt <= 2'h0; // @[FFTDesigns.scala 2131:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FFT_sr_v2_streaming_nrv(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_ready,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
`endif // RANDOMIZE_REG_INIT
  wire  DFT_r_v2_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_1_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_1_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_2_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_2_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_3_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_3_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_4_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_4_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_5_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_5_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_6_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_6_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_7_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_7_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_8_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_8_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_9_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_9_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_10_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_10_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_11_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_11_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_12_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_12_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_13_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_13_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_14_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_14_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_15_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_15_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_16_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_16_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_17_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_17_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_18_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_18_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_19_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_19_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  PermutationsWithStreaming_clock; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_reset; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_0_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_0_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_1_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_1_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_2_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_2_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_3_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_3_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_4_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_4_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_5_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_5_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_6_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_6_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_7_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_7_Im; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_0; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_1; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_2; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_3; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_4; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_5; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_6; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_7; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_8; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_0_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_0_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_1_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_1_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_2_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_2_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_3_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_3_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_4_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_4_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_5_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_5_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_6_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_6_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_7_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_7_Im; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_1_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_5; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_6; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_7; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_8; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_5; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_6; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_7; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_8; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_5; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_6; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_7; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_8; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_5; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_6; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_7; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_8; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_5; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_6; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_7; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_8; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire  TwiddleFactorsStreamed_clock; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_reset; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_7_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_io_in_en_0; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_io_in_en_1; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_7_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_1_clock; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_1_reset; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_7_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_1_io_in_en_0; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_1_io_in_en_1; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_7_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_2_clock; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_2_reset; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_7_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_2_io_in_en_0; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_2_io_in_en_1; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_7_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_3_clock; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_3_reset; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_7_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_3_io_in_en_0; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_3_io_in_en_1; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_7_Im; // @[FFTDesigns.scala 5115:28]
  reg  DFT_regdelays_0_0; // @[FFTDesigns.scala 5094:32]
  reg  DFT_regdelays_1_0; // @[FFTDesigns.scala 5094:32]
  reg  DFT_regdelays_2_0; // @[FFTDesigns.scala 5094:32]
  reg  DFT_regdelays_3_0; // @[FFTDesigns.scala 5094:32]
  reg  DFT_regdelays_4_0; // @[FFTDesigns.scala 5094:32]
  reg  Twid_regdelays_0_0; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_0_1; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_1_0; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_1_1; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_2_0; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_2_1; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_3_0; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_3_1; // @[FFTDesigns.scala 5095:33]
  reg  Perm_regdelays_0_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_4; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_5; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_6; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_7; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_4; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_5; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_6; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_7; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_4; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_5; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_6; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_7; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_4; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_5; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_6; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_7; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_4; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_5; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_6; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_7; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_4; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_5; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_6; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_7; // @[FFTDesigns.scala 5096:33]
  DFT_r_v2 DFT_r_v2 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_clock),
    .reset(DFT_r_v2_reset),
    .io_in_0_Re(DFT_r_v2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_1 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_1_clock),
    .reset(DFT_r_v2_1_reset),
    .io_in_0_Re(DFT_r_v2_1_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_1_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_1_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_1_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_1_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_1_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_1_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_1_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_2 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_2_clock),
    .reset(DFT_r_v2_2_reset),
    .io_in_0_Re(DFT_r_v2_2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_2_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_2_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_3 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_3_clock),
    .reset(DFT_r_v2_3_reset),
    .io_in_0_Re(DFT_r_v2_3_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_3_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_3_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_3_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_3_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_3_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_3_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_3_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_4 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_4_clock),
    .reset(DFT_r_v2_4_reset),
    .io_in_0_Re(DFT_r_v2_4_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_4_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_4_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_4_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_4_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_4_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_4_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_4_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_5 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_5_clock),
    .reset(DFT_r_v2_5_reset),
    .io_in_0_Re(DFT_r_v2_5_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_5_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_5_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_5_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_5_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_5_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_5_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_5_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_6 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_6_clock),
    .reset(DFT_r_v2_6_reset),
    .io_in_0_Re(DFT_r_v2_6_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_6_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_6_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_6_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_6_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_6_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_6_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_6_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_7 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_7_clock),
    .reset(DFT_r_v2_7_reset),
    .io_in_0_Re(DFT_r_v2_7_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_7_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_7_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_7_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_7_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_7_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_7_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_7_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_8 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_8_clock),
    .reset(DFT_r_v2_8_reset),
    .io_in_0_Re(DFT_r_v2_8_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_8_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_8_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_8_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_8_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_8_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_8_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_8_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_9 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_9_clock),
    .reset(DFT_r_v2_9_reset),
    .io_in_0_Re(DFT_r_v2_9_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_9_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_9_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_9_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_9_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_9_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_9_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_9_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_10 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_10_clock),
    .reset(DFT_r_v2_10_reset),
    .io_in_0_Re(DFT_r_v2_10_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_10_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_10_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_10_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_10_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_10_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_10_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_10_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_11 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_11_clock),
    .reset(DFT_r_v2_11_reset),
    .io_in_0_Re(DFT_r_v2_11_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_11_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_11_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_11_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_11_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_11_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_11_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_11_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_12 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_12_clock),
    .reset(DFT_r_v2_12_reset),
    .io_in_0_Re(DFT_r_v2_12_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_12_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_12_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_12_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_12_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_12_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_12_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_12_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_13 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_13_clock),
    .reset(DFT_r_v2_13_reset),
    .io_in_0_Re(DFT_r_v2_13_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_13_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_13_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_13_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_13_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_13_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_13_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_13_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_14 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_14_clock),
    .reset(DFT_r_v2_14_reset),
    .io_in_0_Re(DFT_r_v2_14_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_14_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_14_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_14_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_14_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_14_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_14_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_14_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_15 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_15_clock),
    .reset(DFT_r_v2_15_reset),
    .io_in_0_Re(DFT_r_v2_15_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_15_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_15_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_15_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_15_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_15_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_15_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_15_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_16 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_16_clock),
    .reset(DFT_r_v2_16_reset),
    .io_in_0_Re(DFT_r_v2_16_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_16_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_16_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_16_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_16_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_16_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_16_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_16_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_17 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_17_clock),
    .reset(DFT_r_v2_17_reset),
    .io_in_0_Re(DFT_r_v2_17_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_17_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_17_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_17_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_17_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_17_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_17_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_17_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_18 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_18_clock),
    .reset(DFT_r_v2_18_reset),
    .io_in_0_Re(DFT_r_v2_18_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_18_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_18_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_18_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_18_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_18_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_18_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_18_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_19 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_19_clock),
    .reset(DFT_r_v2_19_reset),
    .io_in_0_Re(DFT_r_v2_19_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_19_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_19_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_19_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_19_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_19_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_19_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_19_io_out_1_Im)
  );
  PermutationsWithStreaming PermutationsWithStreaming ( // @[FFTDesigns.scala 5107:30]
    .clock(PermutationsWithStreaming_clock),
    .reset(PermutationsWithStreaming_reset),
    .io_in_0_Re(PermutationsWithStreaming_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_io_in_7_Im),
    .io_in_en_0(PermutationsWithStreaming_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_io_in_en_8),
    .io_out_0_Re(PermutationsWithStreaming_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_io_out_7_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_1 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_1_clock),
    .reset(PermutationsWithStreaming_1_reset),
    .io_in_0_Re(PermutationsWithStreaming_1_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_1_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_1_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_1_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_1_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_1_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_1_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_1_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_1_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_1_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_1_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_1_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_1_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_1_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_1_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_1_io_in_7_Im),
    .io_in_en_0(PermutationsWithStreaming_1_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_1_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_1_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_1_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_1_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_1_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_1_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_1_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_1_io_in_en_8),
    .io_out_0_Re(PermutationsWithStreaming_1_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_1_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_1_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_1_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_1_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_1_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_1_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_1_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_1_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_1_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_1_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_1_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_1_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_1_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_1_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_1_io_out_7_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_2 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_2_clock),
    .reset(PermutationsWithStreaming_2_reset),
    .io_in_0_Re(PermutationsWithStreaming_2_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_2_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_2_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_2_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_2_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_2_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_2_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_2_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_2_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_2_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_2_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_2_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_2_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_2_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_2_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_2_io_in_7_Im),
    .io_in_en_0(PermutationsWithStreaming_2_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_2_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_2_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_2_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_2_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_2_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_2_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_2_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_2_io_in_en_8),
    .io_out_0_Re(PermutationsWithStreaming_2_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_2_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_2_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_2_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_2_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_2_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_2_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_2_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_2_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_2_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_2_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_2_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_2_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_2_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_2_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_2_io_out_7_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_3 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_3_clock),
    .reset(PermutationsWithStreaming_3_reset),
    .io_in_0_Re(PermutationsWithStreaming_3_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_3_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_3_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_3_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_3_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_3_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_3_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_3_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_3_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_3_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_3_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_3_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_3_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_3_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_3_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_3_io_in_7_Im),
    .io_in_en_0(PermutationsWithStreaming_3_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_3_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_3_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_3_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_3_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_3_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_3_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_3_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_3_io_in_en_8),
    .io_out_0_Re(PermutationsWithStreaming_3_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_3_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_3_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_3_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_3_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_3_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_3_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_3_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_3_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_3_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_3_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_3_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_3_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_3_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_3_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_3_io_out_7_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_4 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_4_clock),
    .reset(PermutationsWithStreaming_4_reset),
    .io_in_0_Re(PermutationsWithStreaming_4_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_4_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_4_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_4_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_4_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_4_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_4_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_4_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_4_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_4_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_4_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_4_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_4_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_4_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_4_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_4_io_in_7_Im),
    .io_in_en_0(PermutationsWithStreaming_4_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_4_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_4_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_4_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_4_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_4_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_4_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_4_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_4_io_in_en_8),
    .io_out_0_Re(PermutationsWithStreaming_4_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_4_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_4_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_4_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_4_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_4_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_4_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_4_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_4_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_4_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_4_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_4_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_4_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_4_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_4_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_4_io_out_7_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_5 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_5_clock),
    .reset(PermutationsWithStreaming_5_reset),
    .io_in_0_Re(PermutationsWithStreaming_5_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_5_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_5_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_5_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_5_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_5_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_5_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_5_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_5_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_5_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_5_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_5_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_5_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_5_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_5_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_5_io_in_7_Im),
    .io_in_en_0(PermutationsWithStreaming_5_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_5_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_5_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_5_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_5_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_5_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_5_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_5_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_5_io_in_en_8),
    .io_out_0_Re(PermutationsWithStreaming_5_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_5_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_5_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_5_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_5_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_5_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_5_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_5_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_5_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_5_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_5_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_5_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_5_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_5_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_5_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_5_io_out_7_Im)
  );
  TwiddleFactorsStreamed TwiddleFactorsStreamed ( // @[FFTDesigns.scala 5115:28]
    .clock(TwiddleFactorsStreamed_clock),
    .reset(TwiddleFactorsStreamed_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_io_in_7_Im),
    .io_in_en_0(TwiddleFactorsStreamed_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_io_out_7_Im)
  );
  TwiddleFactorsStreamed_1 TwiddleFactorsStreamed_1 ( // @[FFTDesigns.scala 5115:28]
    .clock(TwiddleFactorsStreamed_1_clock),
    .reset(TwiddleFactorsStreamed_1_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_1_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_1_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_1_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_1_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_1_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_1_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_1_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_1_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_1_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_1_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_1_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_1_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_1_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_1_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_1_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_1_io_in_7_Im),
    .io_in_en_0(TwiddleFactorsStreamed_1_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_1_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_1_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_1_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_1_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_1_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_1_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_1_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_1_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_1_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_1_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_1_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_1_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_1_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_1_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_1_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_1_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_1_io_out_7_Im)
  );
  TwiddleFactorsStreamed_2 TwiddleFactorsStreamed_2 ( // @[FFTDesigns.scala 5115:28]
    .clock(TwiddleFactorsStreamed_2_clock),
    .reset(TwiddleFactorsStreamed_2_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_2_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_2_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_2_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_2_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_2_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_2_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_2_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_2_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_2_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_2_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_2_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_2_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_2_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_2_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_2_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_2_io_in_7_Im),
    .io_in_en_0(TwiddleFactorsStreamed_2_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_2_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_2_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_2_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_2_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_2_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_2_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_2_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_2_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_2_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_2_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_2_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_2_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_2_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_2_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_2_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_2_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_2_io_out_7_Im)
  );
  TwiddleFactorsStreamed_3 TwiddleFactorsStreamed_3 ( // @[FFTDesigns.scala 5115:28]
    .clock(TwiddleFactorsStreamed_3_clock),
    .reset(TwiddleFactorsStreamed_3_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_3_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_3_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_3_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_3_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_3_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_3_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_3_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_3_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_3_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_3_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_3_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_3_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_3_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_3_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_3_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_3_io_in_7_Im),
    .io_in_en_0(TwiddleFactorsStreamed_3_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_3_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_3_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_3_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_3_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_3_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_3_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_3_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_3_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_3_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_3_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_3_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_3_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_3_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_3_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_3_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_3_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_3_io_out_7_Im)
  );
  assign io_out_0_Re = PermutationsWithStreaming_5_io_out_0_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_0_Im = PermutationsWithStreaming_5_io_out_0_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_1_Re = PermutationsWithStreaming_5_io_out_1_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_1_Im = PermutationsWithStreaming_5_io_out_1_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_2_Re = PermutationsWithStreaming_5_io_out_2_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_2_Im = PermutationsWithStreaming_5_io_out_2_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_3_Re = PermutationsWithStreaming_5_io_out_3_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_3_Im = PermutationsWithStreaming_5_io_out_3_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_4_Re = PermutationsWithStreaming_5_io_out_4_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_4_Im = PermutationsWithStreaming_5_io_out_4_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_5_Re = PermutationsWithStreaming_5_io_out_5_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_5_Im = PermutationsWithStreaming_5_io_out_5_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_6_Re = PermutationsWithStreaming_5_io_out_6_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_6_Im = PermutationsWithStreaming_5_io_out_6_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_7_Re = PermutationsWithStreaming_5_io_out_7_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_7_Im = PermutationsWithStreaming_5_io_out_7_Im; // @[FFTDesigns.scala 5201:12]
  assign DFT_r_v2_clock = clock;
  assign DFT_r_v2_reset = reset;
  assign DFT_r_v2_io_in_0_Re = PermutationsWithStreaming_io_out_0_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_io_in_0_Im = PermutationsWithStreaming_io_out_0_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_io_in_1_Re = PermutationsWithStreaming_io_out_1_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_io_in_1_Im = PermutationsWithStreaming_io_out_1_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_1_clock = clock;
  assign DFT_r_v2_1_reset = reset;
  assign DFT_r_v2_1_io_in_0_Re = PermutationsWithStreaming_io_out_2_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_1_io_in_0_Im = PermutationsWithStreaming_io_out_2_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_1_io_in_1_Re = PermutationsWithStreaming_io_out_3_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_1_io_in_1_Im = PermutationsWithStreaming_io_out_3_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_2_clock = clock;
  assign DFT_r_v2_2_reset = reset;
  assign DFT_r_v2_2_io_in_0_Re = PermutationsWithStreaming_io_out_4_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_2_io_in_0_Im = PermutationsWithStreaming_io_out_4_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_2_io_in_1_Re = PermutationsWithStreaming_io_out_5_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_2_io_in_1_Im = PermutationsWithStreaming_io_out_5_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_3_clock = clock;
  assign DFT_r_v2_3_reset = reset;
  assign DFT_r_v2_3_io_in_0_Re = PermutationsWithStreaming_io_out_6_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_3_io_in_0_Im = PermutationsWithStreaming_io_out_6_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_3_io_in_1_Re = PermutationsWithStreaming_io_out_7_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_3_io_in_1_Im = PermutationsWithStreaming_io_out_7_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_4_clock = clock;
  assign DFT_r_v2_4_reset = reset;
  assign DFT_r_v2_4_io_in_0_Re = TwiddleFactorsStreamed_io_out_0_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_4_io_in_0_Im = TwiddleFactorsStreamed_io_out_0_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_4_io_in_1_Re = TwiddleFactorsStreamed_io_out_1_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_4_io_in_1_Im = TwiddleFactorsStreamed_io_out_1_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_5_clock = clock;
  assign DFT_r_v2_5_reset = reset;
  assign DFT_r_v2_5_io_in_0_Re = TwiddleFactorsStreamed_io_out_2_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_5_io_in_0_Im = TwiddleFactorsStreamed_io_out_2_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_5_io_in_1_Re = TwiddleFactorsStreamed_io_out_3_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_5_io_in_1_Im = TwiddleFactorsStreamed_io_out_3_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_6_clock = clock;
  assign DFT_r_v2_6_reset = reset;
  assign DFT_r_v2_6_io_in_0_Re = TwiddleFactorsStreamed_io_out_4_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_6_io_in_0_Im = TwiddleFactorsStreamed_io_out_4_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_6_io_in_1_Re = TwiddleFactorsStreamed_io_out_5_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_6_io_in_1_Im = TwiddleFactorsStreamed_io_out_5_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_7_clock = clock;
  assign DFT_r_v2_7_reset = reset;
  assign DFT_r_v2_7_io_in_0_Re = TwiddleFactorsStreamed_io_out_6_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_7_io_in_0_Im = TwiddleFactorsStreamed_io_out_6_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_7_io_in_1_Re = TwiddleFactorsStreamed_io_out_7_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_7_io_in_1_Im = TwiddleFactorsStreamed_io_out_7_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_8_clock = clock;
  assign DFT_r_v2_8_reset = reset;
  assign DFT_r_v2_8_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_0_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_8_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_0_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_8_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_1_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_8_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_1_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_9_clock = clock;
  assign DFT_r_v2_9_reset = reset;
  assign DFT_r_v2_9_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_2_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_9_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_2_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_9_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_3_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_9_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_3_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_10_clock = clock;
  assign DFT_r_v2_10_reset = reset;
  assign DFT_r_v2_10_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_4_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_10_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_4_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_10_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_5_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_10_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_5_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_11_clock = clock;
  assign DFT_r_v2_11_reset = reset;
  assign DFT_r_v2_11_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_6_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_11_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_6_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_11_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_7_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_11_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_7_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_12_clock = clock;
  assign DFT_r_v2_12_reset = reset;
  assign DFT_r_v2_12_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_0_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_12_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_0_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_12_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_1_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_12_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_1_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_13_clock = clock;
  assign DFT_r_v2_13_reset = reset;
  assign DFT_r_v2_13_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_2_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_13_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_2_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_13_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_3_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_13_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_3_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_14_clock = clock;
  assign DFT_r_v2_14_reset = reset;
  assign DFT_r_v2_14_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_4_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_14_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_4_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_14_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_5_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_14_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_5_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_15_clock = clock;
  assign DFT_r_v2_15_reset = reset;
  assign DFT_r_v2_15_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_6_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_15_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_6_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_15_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_7_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_15_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_7_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_16_clock = clock;
  assign DFT_r_v2_16_reset = reset;
  assign DFT_r_v2_16_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_0_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_16_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_0_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_16_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_1_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_16_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_1_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_17_clock = clock;
  assign DFT_r_v2_17_reset = reset;
  assign DFT_r_v2_17_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_2_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_17_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_2_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_17_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_3_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_17_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_3_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_18_clock = clock;
  assign DFT_r_v2_18_reset = reset;
  assign DFT_r_v2_18_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_4_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_18_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_4_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_18_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_5_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_18_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_5_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_19_clock = clock;
  assign DFT_r_v2_19_reset = reset;
  assign DFT_r_v2_19_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_6_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_19_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_6_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_19_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_7_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_19_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_7_Im; // @[FFTDesigns.scala 5163:41]
  assign PermutationsWithStreaming_clock = clock;
  assign PermutationsWithStreaming_reset = reset;
  assign PermutationsWithStreaming_io_in_0_Re = io_in_ready ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_0_Im = io_in_ready ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_1_Re = io_in_ready ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_1_Im = io_in_ready ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_2_Re = io_in_ready ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_2_Im = io_in_ready ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_3_Re = io_in_ready ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_3_Im = io_in_ready ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_4_Re = io_in_ready ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_4_Im = io_in_ready ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_5_Re = io_in_ready ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_5_Im = io_in_ready ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_6_Re = io_in_ready ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_6_Im = io_in_ready ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_7_Re = io_in_ready ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_7_Im = io_in_ready ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_en_0 = io_in_ready; // @[FFTDesigns.scala 5123:38]
  assign PermutationsWithStreaming_io_in_en_1 = Perm_regdelays_0_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_2 = Perm_regdelays_0_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_3 = Perm_regdelays_0_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_4 = Perm_regdelays_0_3; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_5 = Perm_regdelays_0_4; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_6 = Perm_regdelays_0_5; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_7 = Perm_regdelays_0_6; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_8 = Perm_regdelays_0_7; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_1_clock = clock;
  assign PermutationsWithStreaming_1_reset = reset;
  assign PermutationsWithStreaming_1_io_in_0_Re = DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_0_Im = DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_1_Re = DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_1_Im = DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_2_Re = DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_2_Im = DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_3_Re = DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_3_Im = DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_4_Re = DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_4_Im = DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_5_Re = DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_5_Im = DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_6_Re = DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_6_Im = DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_7_Re = DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_7_Im = DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_en_0 = DFT_regdelays_0_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_1_io_in_en_1 = Perm_regdelays_1_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_2 = Perm_regdelays_1_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_3 = Perm_regdelays_1_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_4 = Perm_regdelays_1_3; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_5 = Perm_regdelays_1_4; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_6 = Perm_regdelays_1_5; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_7 = Perm_regdelays_1_6; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_8 = Perm_regdelays_1_7; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_2_clock = clock;
  assign PermutationsWithStreaming_2_reset = reset;
  assign PermutationsWithStreaming_2_io_in_0_Re = DFT_r_v2_4_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_0_Im = DFT_r_v2_4_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_1_Re = DFT_r_v2_4_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_1_Im = DFT_r_v2_4_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_2_Re = DFT_r_v2_5_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_2_Im = DFT_r_v2_5_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_3_Re = DFT_r_v2_5_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_3_Im = DFT_r_v2_5_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_4_Re = DFT_r_v2_6_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_4_Im = DFT_r_v2_6_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_5_Re = DFT_r_v2_6_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_5_Im = DFT_r_v2_6_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_6_Re = DFT_r_v2_7_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_6_Im = DFT_r_v2_7_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_7_Re = DFT_r_v2_7_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_7_Im = DFT_r_v2_7_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_en_0 = DFT_regdelays_1_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_2_io_in_en_1 = Perm_regdelays_2_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_2 = Perm_regdelays_2_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_3 = Perm_regdelays_2_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_4 = Perm_regdelays_2_3; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_5 = Perm_regdelays_2_4; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_6 = Perm_regdelays_2_5; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_7 = Perm_regdelays_2_6; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_8 = Perm_regdelays_2_7; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_3_clock = clock;
  assign PermutationsWithStreaming_3_reset = reset;
  assign PermutationsWithStreaming_3_io_in_0_Re = DFT_r_v2_8_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_0_Im = DFT_r_v2_8_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_1_Re = DFT_r_v2_8_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_1_Im = DFT_r_v2_8_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_2_Re = DFT_r_v2_9_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_2_Im = DFT_r_v2_9_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_3_Re = DFT_r_v2_9_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_3_Im = DFT_r_v2_9_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_4_Re = DFT_r_v2_10_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_4_Im = DFT_r_v2_10_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_5_Re = DFT_r_v2_10_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_5_Im = DFT_r_v2_10_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_6_Re = DFT_r_v2_11_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_6_Im = DFT_r_v2_11_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_7_Re = DFT_r_v2_11_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_7_Im = DFT_r_v2_11_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_en_0 = DFT_regdelays_2_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_3_io_in_en_1 = Perm_regdelays_3_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_2 = Perm_regdelays_3_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_3 = Perm_regdelays_3_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_4 = Perm_regdelays_3_3; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_5 = Perm_regdelays_3_4; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_6 = Perm_regdelays_3_5; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_7 = Perm_regdelays_3_6; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_8 = Perm_regdelays_3_7; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_4_clock = clock;
  assign PermutationsWithStreaming_4_reset = reset;
  assign PermutationsWithStreaming_4_io_in_0_Re = DFT_r_v2_12_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_0_Im = DFT_r_v2_12_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_1_Re = DFT_r_v2_12_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_1_Im = DFT_r_v2_12_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_2_Re = DFT_r_v2_13_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_2_Im = DFT_r_v2_13_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_3_Re = DFT_r_v2_13_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_3_Im = DFT_r_v2_13_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_4_Re = DFT_r_v2_14_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_4_Im = DFT_r_v2_14_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_5_Re = DFT_r_v2_14_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_5_Im = DFT_r_v2_14_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_6_Re = DFT_r_v2_15_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_6_Im = DFT_r_v2_15_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_7_Re = DFT_r_v2_15_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_7_Im = DFT_r_v2_15_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_en_0 = DFT_regdelays_3_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_4_io_in_en_1 = Perm_regdelays_4_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_2 = Perm_regdelays_4_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_3 = Perm_regdelays_4_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_4 = Perm_regdelays_4_3; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_5 = Perm_regdelays_4_4; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_6 = Perm_regdelays_4_5; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_7 = Perm_regdelays_4_6; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_8 = Perm_regdelays_4_7; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_5_clock = clock;
  assign PermutationsWithStreaming_5_reset = reset;
  assign PermutationsWithStreaming_5_io_in_0_Re = DFT_r_v2_16_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_0_Im = DFT_r_v2_16_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_1_Re = DFT_r_v2_16_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_1_Im = DFT_r_v2_16_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_2_Re = DFT_r_v2_17_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_2_Im = DFT_r_v2_17_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_3_Re = DFT_r_v2_17_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_3_Im = DFT_r_v2_17_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_4_Re = DFT_r_v2_18_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_4_Im = DFT_r_v2_18_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_5_Re = DFT_r_v2_18_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_5_Im = DFT_r_v2_18_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_6_Re = DFT_r_v2_19_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_6_Im = DFT_r_v2_19_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_7_Re = DFT_r_v2_19_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_7_Im = DFT_r_v2_19_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_en_0 = DFT_regdelays_4_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_5_io_in_en_1 = Perm_regdelays_5_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_2 = Perm_regdelays_5_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_3 = Perm_regdelays_5_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_4 = Perm_regdelays_5_3; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_5 = Perm_regdelays_5_4; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_6 = Perm_regdelays_5_5; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_7 = Perm_regdelays_5_6; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_8 = Perm_regdelays_5_7; // @[FFTDesigns.scala 5144:44]
  assign TwiddleFactorsStreamed_clock = clock;
  assign TwiddleFactorsStreamed_reset = reset;
  assign TwiddleFactorsStreamed_io_in_0_Re = PermutationsWithStreaming_1_io_out_0_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_0_Im = PermutationsWithStreaming_1_io_out_0_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_1_Re = PermutationsWithStreaming_1_io_out_1_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_1_Im = PermutationsWithStreaming_1_io_out_1_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_2_Re = PermutationsWithStreaming_1_io_out_2_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_2_Im = PermutationsWithStreaming_1_io_out_2_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_3_Re = PermutationsWithStreaming_1_io_out_3_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_3_Im = PermutationsWithStreaming_1_io_out_3_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_4_Re = PermutationsWithStreaming_1_io_out_4_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_4_Im = PermutationsWithStreaming_1_io_out_4_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_5_Re = PermutationsWithStreaming_1_io_out_5_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_5_Im = PermutationsWithStreaming_1_io_out_5_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_6_Re = PermutationsWithStreaming_1_io_out_6_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_6_Im = PermutationsWithStreaming_1_io_out_6_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_7_Re = PermutationsWithStreaming_1_io_out_7_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_7_Im = PermutationsWithStreaming_1_io_out_7_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_en_0 = Perm_regdelays_1_7; // @[FFTDesigns.scala 5177:38]
  assign TwiddleFactorsStreamed_io_in_en_1 = Twid_regdelays_0_0; // @[FFTDesigns.scala 5186:36]
  assign TwiddleFactorsStreamed_1_clock = clock;
  assign TwiddleFactorsStreamed_1_reset = reset;
  assign TwiddleFactorsStreamed_1_io_in_0_Re = PermutationsWithStreaming_2_io_out_0_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_0_Im = PermutationsWithStreaming_2_io_out_0_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_1_Re = PermutationsWithStreaming_2_io_out_1_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_1_Im = PermutationsWithStreaming_2_io_out_1_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_2_Re = PermutationsWithStreaming_2_io_out_2_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_2_Im = PermutationsWithStreaming_2_io_out_2_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_3_Re = PermutationsWithStreaming_2_io_out_3_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_3_Im = PermutationsWithStreaming_2_io_out_3_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_4_Re = PermutationsWithStreaming_2_io_out_4_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_4_Im = PermutationsWithStreaming_2_io_out_4_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_5_Re = PermutationsWithStreaming_2_io_out_5_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_5_Im = PermutationsWithStreaming_2_io_out_5_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_6_Re = PermutationsWithStreaming_2_io_out_6_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_6_Im = PermutationsWithStreaming_2_io_out_6_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_7_Re = PermutationsWithStreaming_2_io_out_7_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_7_Im = PermutationsWithStreaming_2_io_out_7_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_en_0 = Perm_regdelays_2_7; // @[FFTDesigns.scala 5181:38]
  assign TwiddleFactorsStreamed_1_io_in_en_1 = Twid_regdelays_1_0; // @[FFTDesigns.scala 5186:36]
  assign TwiddleFactorsStreamed_2_clock = clock;
  assign TwiddleFactorsStreamed_2_reset = reset;
  assign TwiddleFactorsStreamed_2_io_in_0_Re = PermutationsWithStreaming_3_io_out_0_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_0_Im = PermutationsWithStreaming_3_io_out_0_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_1_Re = PermutationsWithStreaming_3_io_out_1_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_1_Im = PermutationsWithStreaming_3_io_out_1_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_2_Re = PermutationsWithStreaming_3_io_out_2_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_2_Im = PermutationsWithStreaming_3_io_out_2_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_3_Re = PermutationsWithStreaming_3_io_out_3_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_3_Im = PermutationsWithStreaming_3_io_out_3_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_4_Re = PermutationsWithStreaming_3_io_out_4_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_4_Im = PermutationsWithStreaming_3_io_out_4_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_5_Re = PermutationsWithStreaming_3_io_out_5_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_5_Im = PermutationsWithStreaming_3_io_out_5_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_6_Re = PermutationsWithStreaming_3_io_out_6_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_6_Im = PermutationsWithStreaming_3_io_out_6_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_7_Re = PermutationsWithStreaming_3_io_out_7_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_7_Im = PermutationsWithStreaming_3_io_out_7_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_en_0 = Perm_regdelays_3_7; // @[FFTDesigns.scala 5181:38]
  assign TwiddleFactorsStreamed_2_io_in_en_1 = Twid_regdelays_2_0; // @[FFTDesigns.scala 5186:36]
  assign TwiddleFactorsStreamed_3_clock = clock;
  assign TwiddleFactorsStreamed_3_reset = reset;
  assign TwiddleFactorsStreamed_3_io_in_0_Re = PermutationsWithStreaming_4_io_out_0_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_0_Im = PermutationsWithStreaming_4_io_out_0_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_1_Re = PermutationsWithStreaming_4_io_out_1_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_1_Im = PermutationsWithStreaming_4_io_out_1_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_2_Re = PermutationsWithStreaming_4_io_out_2_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_2_Im = PermutationsWithStreaming_4_io_out_2_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_3_Re = PermutationsWithStreaming_4_io_out_3_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_3_Im = PermutationsWithStreaming_4_io_out_3_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_4_Re = PermutationsWithStreaming_4_io_out_4_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_4_Im = PermutationsWithStreaming_4_io_out_4_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_5_Re = PermutationsWithStreaming_4_io_out_5_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_5_Im = PermutationsWithStreaming_4_io_out_5_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_6_Re = PermutationsWithStreaming_4_io_out_6_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_6_Im = PermutationsWithStreaming_4_io_out_6_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_7_Re = PermutationsWithStreaming_4_io_out_7_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_7_Im = PermutationsWithStreaming_4_io_out_7_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_en_0 = Perm_regdelays_4_7; // @[FFTDesigns.scala 5181:38]
  assign TwiddleFactorsStreamed_3_io_in_en_1 = Twid_regdelays_3_0; // @[FFTDesigns.scala 5186:36]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_0_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_0_0 <= Perm_regdelays_0_7; // @[FFTDesigns.scala 5153:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_1_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_1_0 <= Twid_regdelays_0_1; // @[FFTDesigns.scala 5160:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_2_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_2_0 <= Twid_regdelays_1_1; // @[FFTDesigns.scala 5160:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_3_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_3_0 <= Twid_regdelays_2_1; // @[FFTDesigns.scala 5160:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_4_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_4_0 <= Twid_regdelays_3_1; // @[FFTDesigns.scala 5160:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_0_0 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_0_0 <= Perm_regdelays_1_7; // @[FFTDesigns.scala 5176:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_0_1 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_0_1 <= Twid_regdelays_0_0; // @[FFTDesigns.scala 5185:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_1_0 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_1_0 <= Perm_regdelays_2_7; // @[FFTDesigns.scala 5180:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_1_1 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_1_1 <= Twid_regdelays_1_0; // @[FFTDesigns.scala 5185:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_2_0 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_2_0 <= Perm_regdelays_3_7; // @[FFTDesigns.scala 5180:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_2_1 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_2_1 <= Twid_regdelays_2_0; // @[FFTDesigns.scala 5185:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_3_0 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_3_0 <= Perm_regdelays_4_7; // @[FFTDesigns.scala 5180:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_3_1 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_3_1 <= Twid_regdelays_3_0; // @[FFTDesigns.scala 5185:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_0 <= io_in_ready; // @[FFTDesigns.scala 5122:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_1 <= Perm_regdelays_0_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_2 <= Perm_regdelays_0_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_3 <= Perm_regdelays_0_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_4 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_4 <= Perm_regdelays_0_3; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_5 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_5 <= Perm_regdelays_0_4; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_6 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_6 <= Perm_regdelays_0_5; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_7 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_7 <= Perm_regdelays_0_6; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_0 <= DFT_regdelays_0_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_1 <= Perm_regdelays_1_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_2 <= Perm_regdelays_1_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_3 <= Perm_regdelays_1_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_4 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_4 <= Perm_regdelays_1_3; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_5 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_5 <= Perm_regdelays_1_4; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_6 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_6 <= Perm_regdelays_1_5; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_7 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_7 <= Perm_regdelays_1_6; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_0 <= DFT_regdelays_1_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_1 <= Perm_regdelays_2_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_2 <= Perm_regdelays_2_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_3 <= Perm_regdelays_2_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_4 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_4 <= Perm_regdelays_2_3; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_5 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_5 <= Perm_regdelays_2_4; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_6 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_6 <= Perm_regdelays_2_5; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_7 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_7 <= Perm_regdelays_2_6; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_0 <= DFT_regdelays_2_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_1 <= Perm_regdelays_3_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_2 <= Perm_regdelays_3_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_3 <= Perm_regdelays_3_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_4 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_4 <= Perm_regdelays_3_3; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_5 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_5 <= Perm_regdelays_3_4; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_6 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_6 <= Perm_regdelays_3_5; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_7 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_7 <= Perm_regdelays_3_6; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_0 <= DFT_regdelays_3_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_1 <= Perm_regdelays_4_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_2 <= Perm_regdelays_4_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_3 <= Perm_regdelays_4_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_4 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_4 <= Perm_regdelays_4_3; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_5 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_5 <= Perm_regdelays_4_4; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_6 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_6 <= Perm_regdelays_4_5; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_7 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_7 <= Perm_regdelays_4_6; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_0 <= DFT_regdelays_4_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_1 <= Perm_regdelays_5_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_2 <= Perm_regdelays_5_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_3 <= Perm_regdelays_5_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_4 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_4 <= Perm_regdelays_5_3; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_5 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_5 <= Perm_regdelays_5_4; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_6 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_6 <= Perm_regdelays_5_5; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_7 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_7 <= Perm_regdelays_5_6; // @[FFTDesigns.scala 5141:32]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DFT_regdelays_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  DFT_regdelays_1_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  DFT_regdelays_2_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  DFT_regdelays_3_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  DFT_regdelays_4_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  Twid_regdelays_0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  Twid_regdelays_0_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  Twid_regdelays_1_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  Twid_regdelays_1_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  Twid_regdelays_2_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  Twid_regdelays_2_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  Twid_regdelays_3_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  Twid_regdelays_3_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  Perm_regdelays_0_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  Perm_regdelays_0_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  Perm_regdelays_0_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  Perm_regdelays_0_3 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  Perm_regdelays_0_4 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  Perm_regdelays_0_5 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  Perm_regdelays_0_6 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  Perm_regdelays_0_7 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  Perm_regdelays_1_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  Perm_regdelays_1_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  Perm_regdelays_1_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  Perm_regdelays_1_3 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  Perm_regdelays_1_4 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  Perm_regdelays_1_5 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  Perm_regdelays_1_6 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  Perm_regdelays_1_7 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  Perm_regdelays_2_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  Perm_regdelays_2_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  Perm_regdelays_2_2 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  Perm_regdelays_2_3 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  Perm_regdelays_2_4 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  Perm_regdelays_2_5 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  Perm_regdelays_2_6 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  Perm_regdelays_2_7 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  Perm_regdelays_3_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  Perm_regdelays_3_1 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  Perm_regdelays_3_2 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  Perm_regdelays_3_3 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  Perm_regdelays_3_4 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  Perm_regdelays_3_5 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  Perm_regdelays_3_6 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  Perm_regdelays_3_7 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  Perm_regdelays_4_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  Perm_regdelays_4_1 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  Perm_regdelays_4_2 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  Perm_regdelays_4_3 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  Perm_regdelays_4_4 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  Perm_regdelays_4_5 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  Perm_regdelays_4_6 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  Perm_regdelays_4_7 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  Perm_regdelays_5_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  Perm_regdelays_5_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  Perm_regdelays_5_2 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  Perm_regdelays_5_3 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  Perm_regdelays_5_4 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  Perm_regdelays_5_5 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  Perm_regdelays_5_6 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  Perm_regdelays_5_7 = _RAND_60[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexSub(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_subber_clock; // @[FPComplex.scala 78:25]
  wire  FP_subber_reset; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 78:25]
  wire  FP_subber_1_clock; // @[FPComplex.scala 78:25]
  wire  FP_subber_1_reset; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_in_a; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_in_b; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_out_s; // @[FPComplex.scala 78:25]
  FP_subber FP_subber ( // @[FPComplex.scala 78:25]
    .clock(FP_subber_clock),
    .reset(FP_subber_reset),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_subber FP_subber_1 ( // @[FPComplex.scala 78:25]
    .clock(FP_subber_1_clock),
    .reset(FP_subber_1_reset),
    .io_in_a(FP_subber_1_io_in_a),
    .io_in_b(FP_subber_1_io_in_b),
    .io_out_s(FP_subber_1_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 85:17]
  assign io_out_s_Im = FP_subber_1_io_out_s; // @[FPComplex.scala 86:17]
  assign FP_subber_clock = clock;
  assign FP_subber_reset = reset;
  assign FP_subber_io_in_a = io_in_a_Re; // @[FPComplex.scala 81:24]
  assign FP_subber_io_in_b = io_in_b_Re; // @[FPComplex.scala 82:24]
  assign FP_subber_1_clock = clock;
  assign FP_subber_1_reset = reset;
  assign FP_subber_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 83:24]
  assign FP_subber_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 84:24]
endmodule
module FPComplexMultiAdder_40(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  assign io_out_Re = io_in_0_Re; // @[FPComplex.scala 521:14]
  assign io_out_Im = io_in_0_Im; // @[FPComplex.scala 521:14]
endmodule
module FPComplexMult_reducable_v2(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 380:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 380:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 380:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 380:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 380:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 380:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 380:33]
  reg [31:0] result_0_Re; // @[FPComplex.scala 391:31]
  reg [31:0] result_0_Im; // @[FPComplex.scala 391:31]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 380:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  assign io_out_s_Re = result_0_Re; // @[FPComplex.scala 400:20]
  assign io_out_s_Im = result_0_Im; // @[FPComplex.scala 400:20]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 381:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 381:24]
  assign cmplx_adj_io_in_adj = 8'h1; // @[FPComplex.scala 384:30]
  assign cmplx_adj_io_is_neg = 1'h1; // @[FPComplex.scala 386:32]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FPComplex.scala 382:29]
  always @(posedge clock) begin
    if (reset) begin // @[FPComplex.scala 391:31]
      result_0_Re <= 32'h0; // @[FPComplex.scala 391:31]
    end else begin
      result_0_Re <= cmplx_adj_io_out_Re; // @[FPComplex.scala 394:25]
    end
    if (reset) begin // @[FPComplex.scala 391:31]
      result_0_Im <= 32'h0; // @[FPComplex.scala 391:31]
    end else begin
      result_0_Im <= cmplx_adj_io_out_Im; // @[FPComplex.scala 394:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  result_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  result_0_Im = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMult_reducable_v2_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 340:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 340:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 340:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 340:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 340:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 340:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 340:33]
  wire  FP_multiplier_clock; // @[FPComplex.scala 368:29]
  wire  FP_multiplier_reset; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 368:29]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 368:29]
  wire  FP_multiplier_1_reset; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 368:29]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 340:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 368:29]
    .clock(FP_multiplier_clock),
    .reset(FP_multiplier_reset),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 368:29]
    .clock(FP_multiplier_1_clock),
    .reset(FP_multiplier_1_reset),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  assign io_out_s_Re = FP_multiplier_io_out_s; // @[FPComplex.scala 375:21]
  assign io_out_s_Im = FP_multiplier_1_io_out_s; // @[FPComplex.scala 376:21]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 341:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 341:24]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FPComplex.scala 365:30]
  assign cmplx_adj_io_is_neg = 1'h0; // @[FPComplex.scala 366:30]
  assign cmplx_adj_io_is_flip = 1'h1; // @[FPComplex.scala 342:29]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_reset = reset;
  assign FP_multiplier_io_in_a = cmplx_adj_io_out_Re; // @[FPComplex.scala 371:29]
  assign FP_multiplier_io_in_b = 32'hbf5db3d6; // @[FPComplex.scala 372:29]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_reset = reset;
  assign FP_multiplier_1_io_in_a = cmplx_adj_io_out_Im; // @[FPComplex.scala 373:29]
  assign FP_multiplier_1_io_in_b = 32'hbf5db3d6; // @[FPComplex.scala 374:29]
endmodule
module DFT_r_v2_20(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  FPComplexAdder_clock; // @[FFTDesigns.scala 258:34]
  wire  FPComplexAdder_reset; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_a_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_a_Im; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_b_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_b_Im; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 258:34]
  wire  FPComplexSub_clock; // @[FFTDesigns.scala 261:34]
  wire  FPComplexSub_reset; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_a_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_a_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_b_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_b_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_out_s_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_out_s_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexMultiAdder_io_in_0_Re; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_in_0_Im; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 275:36]
  wire  FPComplexMult_reducable_v2_clock; // @[FFTDesigns.scala 294:39]
  wire  FPComplexMult_reducable_v2_reset; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Re; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Im; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 294:39]
  wire  FPComplexMult_reducable_v2_1_clock; // @[FFTDesigns.scala 297:39]
  wire  FPComplexMult_reducable_v2_1_reset; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Re; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Im; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 297:39]
  wire  FPComplexAdder_reducable_clock; // @[FFTDesigns.scala 338:34]
  wire  FPComplexAdder_reducable_reset; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_a_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_a_Im; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_b_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_b_Im; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_out_s_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_out_s_Im; // @[FFTDesigns.scala 338:34]
  wire  FPComplexSub_reducable_clock; // @[FFTDesigns.scala 341:34]
  wire  FPComplexSub_reducable_reset; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_a_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_a_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_b_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_b_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_out_s_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_out_s_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_in_0_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_in_0_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_out_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_out_Im; // @[FFTDesigns.scala 394:29]
  wire  FPComplexAdder_1_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_1_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_2_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_2_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_3_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_3_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  reg [31:0] initial_layer_out_0_0_Re; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_0_0_Im; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_1_0_Re; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_1_0_Im; // @[FFTDesigns.scala 276:84]
  reg [31:0] finallayer_0_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_0_Im; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_1_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_1_Im; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_2_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_2_Im; // @[FFTDesigns.scala 421:31]
  FPComplexAdder FPComplexAdder ( // @[FFTDesigns.scala 258:34]
    .clock(FPComplexAdder_clock),
    .reset(FPComplexAdder_reset),
    .io_in_a_Re(FPComplexAdder_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_io_out_s_Im)
  );
  FPComplexSub FPComplexSub ( // @[FFTDesigns.scala 261:34]
    .clock(FPComplexSub_clock),
    .reset(FPComplexSub_reset),
    .io_in_a_Re(FPComplexSub_io_in_a_Re),
    .io_in_a_Im(FPComplexSub_io_in_a_Im),
    .io_in_b_Re(FPComplexSub_io_in_b_Re),
    .io_in_b_Im(FPComplexSub_io_in_b_Im),
    .io_out_s_Re(FPComplexSub_io_out_s_Re),
    .io_out_s_Im(FPComplexSub_io_out_s_Im)
  );
  FPComplexMultiAdder_40 FPComplexMultiAdder ( // @[FFTDesigns.scala 275:36]
    .io_in_0_Re(FPComplexMultiAdder_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_io_out_Im)
  );
  FPComplexMult_reducable_v2 FPComplexMult_reducable_v2 ( // @[FFTDesigns.scala 294:39]
    .clock(FPComplexMult_reducable_v2_clock),
    .reset(FPComplexMult_reducable_v2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_1 FPComplexMult_reducable_v2_1 ( // @[FFTDesigns.scala 297:39]
    .clock(FPComplexMult_reducable_v2_1_clock),
    .reset(FPComplexMult_reducable_v2_1_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_1_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_1_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_reducable ( // @[FFTDesigns.scala 338:34]
    .clock(FPComplexAdder_reducable_clock),
    .reset(FPComplexAdder_reducable_reset),
    .io_in_a_Re(FPComplexAdder_reducable_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_reducable_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_reducable_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_reducable_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_reducable_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_reducable_io_out_s_Im)
  );
  FPComplexSub FPComplexSub_reducable ( // @[FFTDesigns.scala 341:34]
    .clock(FPComplexSub_reducable_clock),
    .reset(FPComplexSub_reducable_reset),
    .io_in_a_Re(FPComplexSub_reducable_io_in_a_Re),
    .io_in_a_Im(FPComplexSub_reducable_io_in_a_Im),
    .io_in_b_Re(FPComplexSub_reducable_io_in_b_Re),
    .io_in_b_Im(FPComplexSub_reducable_io_in_b_Im),
    .io_out_s_Re(FPComplexSub_reducable_io_out_s_Re),
    .io_out_s_Im(FPComplexSub_reducable_io_out_s_Im)
  );
  FPComplexMultiAdder_40 FPComplexMultiAdder_1 ( // @[FFTDesigns.scala 394:29]
    .io_in_0_Re(FPComplexMultiAdder_1_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_1_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_1_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_1_io_out_Im)
  );
  FPComplexMultiAdder_40 FPComplexMultiAdder_2 ( // @[FFTDesigns.scala 394:29]
    .io_in_0_Re(FPComplexMultiAdder_2_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_2_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_2_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_2_io_out_Im)
  );
  FPComplexAdder FPComplexAdder_1 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_1_clock),
    .reset(FPComplexAdder_1_reset),
    .io_in_a_Re(FPComplexAdder_1_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_1_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_1_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_1_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_1_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_1_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_2 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_2_clock),
    .reset(FPComplexAdder_2_reset),
    .io_in_a_Re(FPComplexAdder_2_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_2_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_2_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_2_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_2_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_2_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_3 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_3_clock),
    .reset(FPComplexAdder_3_reset),
    .io_in_a_Re(FPComplexAdder_3_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_3_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_3_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_3_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_3_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_3_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexAdder_1_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_0_Im = FPComplexAdder_1_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign io_out_1_Re = FPComplexAdder_2_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_1_Im = FPComplexAdder_2_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign io_out_2_Re = FPComplexAdder_3_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_2_Im = FPComplexAdder_3_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign FPComplexAdder_clock = clock;
  assign FPComplexAdder_reset = reset;
  assign FPComplexAdder_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 268:38]
  assign FPComplexAdder_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 268:38]
  assign FPComplexAdder_io_in_b_Re = io_in_2_Re; // @[FFTDesigns.scala 269:38]
  assign FPComplexAdder_io_in_b_Im = io_in_2_Im; // @[FFTDesigns.scala 269:38]
  assign FPComplexSub_clock = clock;
  assign FPComplexSub_reset = reset;
  assign FPComplexSub_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 270:38]
  assign FPComplexSub_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 270:38]
  assign FPComplexSub_io_in_b_Re = io_in_2_Re; // @[FFTDesigns.scala 271:38]
  assign FPComplexSub_io_in_b_Im = io_in_2_Im; // @[FFTDesigns.scala 271:38]
  assign FPComplexMultiAdder_io_in_0_Re = initial_layer_out_1_0_Re; // @[FFTDesigns.scala 290:27]
  assign FPComplexMultiAdder_io_in_0_Im = initial_layer_out_1_0_Im; // @[FFTDesigns.scala 290:27]
  assign FPComplexMult_reducable_v2_clock = clock;
  assign FPComplexMult_reducable_v2_reset = reset;
  assign FPComplexMult_reducable_v2_io_in_a_Re = FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 320:34]
  assign FPComplexMult_reducable_v2_io_in_a_Im = FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 320:34]
  assign FPComplexMult_reducable_v2_1_clock = clock;
  assign FPComplexMult_reducable_v2_1_reset = reset;
  assign FPComplexMult_reducable_v2_1_io_in_a_Re = FPComplexSub_io_out_s_Re; // @[FFTDesigns.scala 323:34]
  assign FPComplexMult_reducable_v2_1_io_in_a_Im = FPComplexSub_io_out_s_Im; // @[FFTDesigns.scala 323:34]
  assign FPComplexAdder_reducable_clock = clock;
  assign FPComplexAdder_reducable_reset = reset;
  assign FPComplexAdder_reducable_io_in_a_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 366:36]
  assign FPComplexAdder_reducable_io_in_a_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 366:36]
  assign FPComplexAdder_reducable_io_in_b_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 367:36]
  assign FPComplexAdder_reducable_io_in_b_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 367:36]
  assign FPComplexSub_reducable_clock = clock;
  assign FPComplexSub_reducable_reset = reset;
  assign FPComplexSub_reducable_io_in_a_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 368:36]
  assign FPComplexSub_reducable_io_in_a_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 368:36]
  assign FPComplexSub_reducable_io_in_b_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 369:36]
  assign FPComplexSub_reducable_io_in_b_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 369:36]
  assign FPComplexMultiAdder_1_io_in_0_Re = FPComplexAdder_reducable_io_out_s_Re; // @[FFTDesigns.scala 402:36]
  assign FPComplexMultiAdder_1_io_in_0_Im = FPComplexAdder_reducable_io_out_s_Im; // @[FFTDesigns.scala 402:36]
  assign FPComplexMultiAdder_2_io_in_0_Re = FPComplexSub_reducable_io_out_s_Re; // @[FFTDesigns.scala 404:61]
  assign FPComplexMultiAdder_2_io_in_0_Im = FPComplexSub_reducable_io_out_s_Im; // @[FFTDesigns.scala 404:61]
  assign FPComplexAdder_1_clock = clock;
  assign FPComplexAdder_1_reset = reset;
  assign FPComplexAdder_1_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_1_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_1_io_in_b_Re = FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_1_io_in_b_Im = FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_2_clock = clock;
  assign FPComplexAdder_2_reset = reset;
  assign FPComplexAdder_2_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_2_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_2_io_in_b_Re = FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_2_io_in_b_Im = FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_3_clock = clock;
  assign FPComplexAdder_3_reset = reset;
  assign FPComplexAdder_3_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_3_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_3_io_in_b_Re = FPComplexMultiAdder_2_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_3_io_in_b_Im = FPComplexMultiAdder_2_io_out_Im; // @[FFTDesigns.scala 431:35]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_0_0_Re <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_0_0_Re <= FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 281:37]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_0_0_Im <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_0_0_Im <= FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 281:37]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_1_0_Re <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_1_0_Re <= initial_layer_out_0_0_Re; // @[FFTDesigns.scala 284:32]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_1_0_Im <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_1_0_Im <= initial_layer_out_0_0_Im; // @[FFTDesigns.scala 284:32]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_0_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_0_Re <= io_in_0_Re; // @[FFTDesigns.scala 424:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_0_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_0_Im <= io_in_0_Im; // @[FFTDesigns.scala 424:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_1_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_1_Re <= finallayer_0_Re; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_1_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_1_Im <= finallayer_0_Im; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_2_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_2_Re <= finallayer_1_Re; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_2_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_2_Im <= finallayer_1_Im; // @[FFTDesigns.scala 426:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  initial_layer_out_0_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  initial_layer_out_0_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  initial_layer_out_1_0_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  initial_layer_out_1_0_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  finallayer_0_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  finallayer_0_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  finallayer_1_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  finallayer_1_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  finallayer_2_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  finallayer_2_Im = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_Block_96(
  input         clock,
  input  [4:0]  io_in_raddr,
  input  [4:0]  io_in_waddr,
  input  [31:0] io_in_data_Re,
  input  [31:0] io_in_data_Im,
  input         io_re,
  input         io_wr,
  input         io_en,
  output [31:0] io_out_data_Re,
  output [31:0] io_out_data_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_0_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_8_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_8_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_9_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_9_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_10_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_10_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_11_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_11_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_12_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_12_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_13_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_13_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_14_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_14_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_15_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_15_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_16_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_16_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_17_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_17_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_18_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_18_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_19_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_19_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_20_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_20_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_21_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_21_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_22_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_22_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_23_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_23_Im; // @[FFTDesigns.scala 3286:18]
  wire [31:0] _GEN_97 = 5'h1 == io_in_raddr ? mem_1_Im : mem_0_Im; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_98 = 5'h2 == io_in_raddr ? mem_2_Im : _GEN_97; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_99 = 5'h3 == io_in_raddr ? mem_3_Im : _GEN_98; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_100 = 5'h4 == io_in_raddr ? mem_4_Im : _GEN_99; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_101 = 5'h5 == io_in_raddr ? mem_5_Im : _GEN_100; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_102 = 5'h6 == io_in_raddr ? mem_6_Im : _GEN_101; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_103 = 5'h7 == io_in_raddr ? mem_7_Im : _GEN_102; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_104 = 5'h8 == io_in_raddr ? mem_8_Im : _GEN_103; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_105 = 5'h9 == io_in_raddr ? mem_9_Im : _GEN_104; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_106 = 5'ha == io_in_raddr ? mem_10_Im : _GEN_105; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_107 = 5'hb == io_in_raddr ? mem_11_Im : _GEN_106; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_108 = 5'hc == io_in_raddr ? mem_12_Im : _GEN_107; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_109 = 5'hd == io_in_raddr ? mem_13_Im : _GEN_108; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_110 = 5'he == io_in_raddr ? mem_14_Im : _GEN_109; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_111 = 5'hf == io_in_raddr ? mem_15_Im : _GEN_110; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_112 = 5'h10 == io_in_raddr ? mem_16_Im : _GEN_111; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_113 = 5'h11 == io_in_raddr ? mem_17_Im : _GEN_112; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_114 = 5'h12 == io_in_raddr ? mem_18_Im : _GEN_113; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_115 = 5'h13 == io_in_raddr ? mem_19_Im : _GEN_114; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_116 = 5'h14 == io_in_raddr ? mem_20_Im : _GEN_115; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_117 = 5'h15 == io_in_raddr ? mem_21_Im : _GEN_116; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_118 = 5'h16 == io_in_raddr ? mem_22_Im : _GEN_117; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_119 = 5'h17 == io_in_raddr ? mem_23_Im : _GEN_118; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_121 = 5'h1 == io_in_raddr ? mem_1_Re : mem_0_Re; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_122 = 5'h2 == io_in_raddr ? mem_2_Re : _GEN_121; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_123 = 5'h3 == io_in_raddr ? mem_3_Re : _GEN_122; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_124 = 5'h4 == io_in_raddr ? mem_4_Re : _GEN_123; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_125 = 5'h5 == io_in_raddr ? mem_5_Re : _GEN_124; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_126 = 5'h6 == io_in_raddr ? mem_6_Re : _GEN_125; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_127 = 5'h7 == io_in_raddr ? mem_7_Re : _GEN_126; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_128 = 5'h8 == io_in_raddr ? mem_8_Re : _GEN_127; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_129 = 5'h9 == io_in_raddr ? mem_9_Re : _GEN_128; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_130 = 5'ha == io_in_raddr ? mem_10_Re : _GEN_129; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_131 = 5'hb == io_in_raddr ? mem_11_Re : _GEN_130; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_132 = 5'hc == io_in_raddr ? mem_12_Re : _GEN_131; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_133 = 5'hd == io_in_raddr ? mem_13_Re : _GEN_132; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_134 = 5'he == io_in_raddr ? mem_14_Re : _GEN_133; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_135 = 5'hf == io_in_raddr ? mem_15_Re : _GEN_134; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_136 = 5'h10 == io_in_raddr ? mem_16_Re : _GEN_135; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_137 = 5'h11 == io_in_raddr ? mem_17_Re : _GEN_136; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_138 = 5'h12 == io_in_raddr ? mem_18_Re : _GEN_137; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_139 = 5'h13 == io_in_raddr ? mem_19_Re : _GEN_138; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_140 = 5'h14 == io_in_raddr ? mem_20_Re : _GEN_139; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_141 = 5'h15 == io_in_raddr ? mem_21_Re : _GEN_140; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_142 = 5'h16 == io_in_raddr ? mem_22_Re : _GEN_141; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_143 = 5'h17 == io_in_raddr ? mem_23_Re : _GEN_142; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_144 = io_re ? _GEN_119 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3295:24]
  wire [31:0] _GEN_145 = io_re ? _GEN_143 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3294:24]
  assign io_out_data_Re = io_en ? _GEN_145 : 32'h0; // @[FFTDesigns.scala 3287:16 3298:22]
  assign io_out_data_Im = io_en ? _GEN_144 : 32'h0; // @[FFTDesigns.scala 3287:16 3299:22]
  always @(posedge clock) begin
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h8 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_8_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h8 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_8_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h9 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_9_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h9 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_9_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'ha == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_10_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'ha == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_10_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'hb == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_11_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'hb == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_11_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'hc == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_12_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'hc == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_12_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'hd == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_13_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'hd == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_13_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'he == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_14_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'he == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_14_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'hf == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_15_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'hf == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_15_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h10 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_16_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h10 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_16_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h11 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_17_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h11 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_17_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h12 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_18_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h12 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_18_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h13 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_19_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h13 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_19_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h14 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_20_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h14 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_20_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h15 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_21_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h15 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_21_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h16 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_22_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h16 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_22_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h17 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_23_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (5'h17 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_23_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_3_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_4_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_4_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_5_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_5_Im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_6_Re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_6_Im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_7_Re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_7_Im = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mem_8_Re = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mem_8_Im = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_9_Re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mem_9_Im = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mem_10_Re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mem_10_Im = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_11_Re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mem_11_Im = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  mem_12_Re = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  mem_12_Im = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  mem_13_Re = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mem_13_Im = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mem_14_Re = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mem_14_Im = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mem_15_Re = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mem_15_Im = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mem_16_Re = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mem_16_Im = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mem_17_Re = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mem_17_Im = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mem_18_Re = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mem_18_Im = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mem_19_Re = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mem_19_Im = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mem_20_Re = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mem_20_Im = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mem_21_Re = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mem_21_Im = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mem_22_Re = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mem_22_Im = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mem_23_Re = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mem_23_Im = _RAND_47[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module M0_Config_ROM_6(
  input  [3:0] io_in_cnt,
  output [4:0] io_out_0,
  output [4:0] io_out_1,
  output [4:0] io_out_2,
  output [4:0] io_out_3,
  output [4:0] io_out_4,
  output [4:0] io_out_5,
  output [4:0] io_out_6,
  output [4:0] io_out_7
);
  wire [4:0] _GEN_1 = 4'h1 == io_in_cnt ? 5'h1 : 5'h0; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_2 = 4'h2 == io_in_cnt ? 5'h2 : _GEN_1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_3 = 4'h3 == io_in_cnt ? 5'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_4 = 4'h4 == io_in_cnt ? 5'h4 : _GEN_3; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_5 = 4'h5 == io_in_cnt ? 5'h5 : _GEN_4; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_6 = 4'h6 == io_in_cnt ? 5'h6 : _GEN_5; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_7 = 4'h7 == io_in_cnt ? 5'h7 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_8 = 4'h8 == io_in_cnt ? 5'h8 : _GEN_7; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_9 = 4'h9 == io_in_cnt ? 5'h9 : _GEN_8; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_10 = 4'ha == io_in_cnt ? 5'ha : _GEN_9; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_13 = 4'h1 == io_in_cnt ? 5'h2 : 5'h1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_14 = 4'h2 == io_in_cnt ? 5'h3 : _GEN_13; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_15 = 4'h3 == io_in_cnt ? 5'h4 : _GEN_14; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_16 = 4'h4 == io_in_cnt ? 5'h5 : _GEN_15; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_17 = 4'h5 == io_in_cnt ? 5'h6 : _GEN_16; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_18 = 4'h6 == io_in_cnt ? 5'h7 : _GEN_17; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_19 = 4'h7 == io_in_cnt ? 5'h8 : _GEN_18; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_20 = 4'h8 == io_in_cnt ? 5'h9 : _GEN_19; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_21 = 4'h9 == io_in_cnt ? 5'ha : _GEN_20; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_22 = 4'ha == io_in_cnt ? 5'hb : _GEN_21; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_25 = 4'h1 == io_in_cnt ? 5'h3 : 5'h2; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_26 = 4'h2 == io_in_cnt ? 5'h4 : _GEN_25; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_27 = 4'h3 == io_in_cnt ? 5'h5 : _GEN_26; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_28 = 4'h4 == io_in_cnt ? 5'h6 : _GEN_27; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_29 = 4'h5 == io_in_cnt ? 5'h7 : _GEN_28; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_30 = 4'h6 == io_in_cnt ? 5'h8 : _GEN_29; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_31 = 4'h7 == io_in_cnt ? 5'h9 : _GEN_30; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_32 = 4'h8 == io_in_cnt ? 5'ha : _GEN_31; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_33 = 4'h9 == io_in_cnt ? 5'hb : _GEN_32; // @[FFTDesigns.scala 3227:{17,17}]
  wire [4:0] _GEN_34 = 4'ha == io_in_cnt ? 5'h0 : _GEN_33; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_0 = 4'hb == io_in_cnt ? 5'hb : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_1 = 4'hb == io_in_cnt ? 5'h0 : _GEN_22; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_2 = 4'hb == io_in_cnt ? 5'h1 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_3 = 4'hb == io_in_cnt ? 5'hb : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_4 = 4'hb == io_in_cnt ? 5'h0 : _GEN_22; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_5 = 4'hb == io_in_cnt ? 5'h1 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_6 = 4'hb == io_in_cnt ? 5'hb : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_7 = 4'hb == io_in_cnt ? 5'h0 : _GEN_22; // @[FFTDesigns.scala 3227:{17,17}]
endmodule
module M1_Config_ROM_6(
  input  [3:0] io_in_cnt,
  output [4:0] io_out_0,
  output [4:0] io_out_1,
  output [4:0] io_out_2,
  output [4:0] io_out_3,
  output [4:0] io_out_4,
  output [4:0] io_out_5,
  output [4:0] io_out_6,
  output [4:0] io_out_7
);
  wire [4:0] _GEN_1 = 4'h1 == io_in_cnt ? 5'h9 : 5'h0; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_2 = 4'h2 == io_in_cnt ? 5'h5 : _GEN_1; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_3 = 4'h3 == io_in_cnt ? 5'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_4 = 4'h4 == io_in_cnt ? 5'ha : _GEN_3; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_5 = 4'h5 == io_in_cnt ? 5'h6 : _GEN_4; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_6 = 4'h6 == io_in_cnt ? 5'h2 : _GEN_5; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_7 = 4'h7 == io_in_cnt ? 5'hb : _GEN_6; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_8 = 4'h8 == io_in_cnt ? 5'h7 : _GEN_7; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_9 = 4'h9 == io_in_cnt ? 5'h3 : _GEN_8; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_10 = 4'ha == io_in_cnt ? 5'h8 : _GEN_9; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_25 = 4'h1 == io_in_cnt ? 5'h8 : 5'h0; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_26 = 4'h2 == io_in_cnt ? 5'h5 : _GEN_25; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_27 = 4'h3 == io_in_cnt ? 5'h1 : _GEN_26; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_28 = 4'h4 == io_in_cnt ? 5'h9 : _GEN_27; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_29 = 4'h5 == io_in_cnt ? 5'h6 : _GEN_28; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_30 = 4'h6 == io_in_cnt ? 5'h2 : _GEN_29; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_31 = 4'h7 == io_in_cnt ? 5'ha : _GEN_30; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_32 = 4'h8 == io_in_cnt ? 5'h7 : _GEN_31; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_33 = 4'h9 == io_in_cnt ? 5'h3 : _GEN_32; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_34 = 4'ha == io_in_cnt ? 5'hb : _GEN_33; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_62 = 4'h2 == io_in_cnt ? 5'h4 : _GEN_25; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_63 = 4'h3 == io_in_cnt ? 5'h1 : _GEN_62; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_64 = 4'h4 == io_in_cnt ? 5'h9 : _GEN_63; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_65 = 4'h5 == io_in_cnt ? 5'h5 : _GEN_64; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_66 = 4'h6 == io_in_cnt ? 5'h2 : _GEN_65; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_67 = 4'h7 == io_in_cnt ? 5'ha : _GEN_66; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_68 = 4'h8 == io_in_cnt ? 5'h6 : _GEN_67; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_69 = 4'h9 == io_in_cnt ? 5'h3 : _GEN_68; // @[FFTDesigns.scala 3250:{17,17}]
  wire [4:0] _GEN_70 = 4'ha == io_in_cnt ? 5'hb : _GEN_69; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_0 = 4'hb == io_in_cnt ? 5'h4 : _GEN_10; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_1 = 4'hb == io_in_cnt ? 5'h4 : _GEN_10; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_2 = 4'hb == io_in_cnt ? 5'h4 : _GEN_34; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_3 = 4'hb == io_in_cnt ? 5'h4 : _GEN_34; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_4 = 4'hb == io_in_cnt ? 5'h4 : _GEN_34; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_5 = 4'hb == io_in_cnt ? 5'h7 : _GEN_70; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_6 = 4'hb == io_in_cnt ? 5'h7 : _GEN_70; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_7 = 4'hb == io_in_cnt ? 5'h7 : _GEN_70; // @[FFTDesigns.scala 3250:{17,17}]
endmodule
module Streaming_Permute_Config_6(
  input  [3:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6
);
  wire [2:0] _GEN_1 = 4'h1 == io_in_cnt ? 3'h2 : 3'h0; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_2 = 4'h2 == io_in_cnt ? 3'h5 : _GEN_1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_3 = 4'h3 == io_in_cnt ? 3'h0 : _GEN_2; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_4 = 4'h4 == io_in_cnt ? 3'h2 : _GEN_3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_5 = 4'h5 == io_in_cnt ? 3'h5 : _GEN_4; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_6 = 4'h6 == io_in_cnt ? 3'h0 : _GEN_5; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_7 = 4'h7 == io_in_cnt ? 3'h2 : _GEN_6; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_8 = 4'h8 == io_in_cnt ? 3'h5 : _GEN_7; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_9 = 4'h9 == io_in_cnt ? 3'h0 : _GEN_8; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_10 = 4'ha == io_in_cnt ? 3'h2 : _GEN_9; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_13 = 4'h1 == io_in_cnt ? 3'h5 : 3'h3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_14 = 4'h2 == io_in_cnt ? 3'h0 : _GEN_13; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_15 = 4'h3 == io_in_cnt ? 3'h3 : _GEN_14; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_16 = 4'h4 == io_in_cnt ? 3'h5 : _GEN_15; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_17 = 4'h5 == io_in_cnt ? 3'h0 : _GEN_16; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_18 = 4'h6 == io_in_cnt ? 3'h3 : _GEN_17; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_19 = 4'h7 == io_in_cnt ? 3'h5 : _GEN_18; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_20 = 4'h8 == io_in_cnt ? 3'h0 : _GEN_19; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_21 = 4'h9 == io_in_cnt ? 3'h3 : _GEN_20; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_22 = 4'ha == io_in_cnt ? 3'h5 : _GEN_21; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_25 = 4'h1 == io_in_cnt ? 3'h0 : 3'h6; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_26 = 4'h2 == io_in_cnt ? 3'h3 : _GEN_25; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_27 = 4'h3 == io_in_cnt ? 3'h6 : _GEN_26; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_28 = 4'h4 == io_in_cnt ? 3'h0 : _GEN_27; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_29 = 4'h5 == io_in_cnt ? 3'h3 : _GEN_28; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_30 = 4'h6 == io_in_cnt ? 3'h6 : _GEN_29; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_31 = 4'h7 == io_in_cnt ? 3'h0 : _GEN_30; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_32 = 4'h8 == io_in_cnt ? 3'h3 : _GEN_31; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_33 = 4'h9 == io_in_cnt ? 3'h6 : _GEN_32; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_34 = 4'ha == io_in_cnt ? 3'h0 : _GEN_33; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_37 = 4'h1 == io_in_cnt ? 3'h3 : 3'h1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_38 = 4'h2 == io_in_cnt ? 3'h6 : _GEN_37; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_39 = 4'h3 == io_in_cnt ? 3'h1 : _GEN_38; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_40 = 4'h4 == io_in_cnt ? 3'h3 : _GEN_39; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_41 = 4'h5 == io_in_cnt ? 3'h6 : _GEN_40; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_42 = 4'h6 == io_in_cnt ? 3'h1 : _GEN_41; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_43 = 4'h7 == io_in_cnt ? 3'h3 : _GEN_42; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_44 = 4'h8 == io_in_cnt ? 3'h6 : _GEN_43; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_45 = 4'h9 == io_in_cnt ? 3'h1 : _GEN_44; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_46 = 4'ha == io_in_cnt ? 3'h3 : _GEN_45; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_49 = 4'h1 == io_in_cnt ? 3'h6 : 3'h4; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_50 = 4'h2 == io_in_cnt ? 3'h1 : _GEN_49; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_51 = 4'h3 == io_in_cnt ? 3'h4 : _GEN_50; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_52 = 4'h4 == io_in_cnt ? 3'h6 : _GEN_51; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_53 = 4'h5 == io_in_cnt ? 3'h1 : _GEN_52; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_54 = 4'h6 == io_in_cnt ? 3'h4 : _GEN_53; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_55 = 4'h7 == io_in_cnt ? 3'h6 : _GEN_54; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_56 = 4'h8 == io_in_cnt ? 3'h1 : _GEN_55; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_57 = 4'h9 == io_in_cnt ? 3'h4 : _GEN_56; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_58 = 4'ha == io_in_cnt ? 3'h6 : _GEN_57; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_61 = 4'h1 == io_in_cnt ? 3'h1 : 3'h7; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_62 = 4'h2 == io_in_cnt ? 3'h4 : _GEN_61; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_63 = 4'h3 == io_in_cnt ? 3'h7 : _GEN_62; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_64 = 4'h4 == io_in_cnt ? 3'h1 : _GEN_63; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_65 = 4'h5 == io_in_cnt ? 3'h4 : _GEN_64; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_66 = 4'h6 == io_in_cnt ? 3'h7 : _GEN_65; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_67 = 4'h7 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_68 = 4'h8 == io_in_cnt ? 3'h4 : _GEN_67; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_69 = 4'h9 == io_in_cnt ? 3'h7 : _GEN_68; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_70 = 4'ha == io_in_cnt ? 3'h1 : _GEN_69; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_73 = 4'h1 == io_in_cnt ? 3'h4 : 3'h2; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_74 = 4'h2 == io_in_cnt ? 3'h7 : _GEN_73; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_75 = 4'h3 == io_in_cnt ? 3'h2 : _GEN_74; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_76 = 4'h4 == io_in_cnt ? 3'h4 : _GEN_75; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_77 = 4'h5 == io_in_cnt ? 3'h7 : _GEN_76; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_78 = 4'h6 == io_in_cnt ? 3'h2 : _GEN_77; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_79 = 4'h7 == io_in_cnt ? 3'h4 : _GEN_78; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_80 = 4'h8 == io_in_cnt ? 3'h7 : _GEN_79; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_81 = 4'h9 == io_in_cnt ? 3'h2 : _GEN_80; // @[FFTDesigns.scala 3273:{17,17}]
  wire [2:0] _GEN_82 = 4'ha == io_in_cnt ? 3'h4 : _GEN_81; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_0 = 4'hb == io_in_cnt ? 3'h5 : _GEN_10; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_1 = 4'hb == io_in_cnt ? 3'h0 : _GEN_22; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_2 = 4'hb == io_in_cnt ? 3'h3 : _GEN_34; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_3 = 4'hb == io_in_cnt ? 3'h6 : _GEN_46; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_4 = 4'hb == io_in_cnt ? 3'h1 : _GEN_58; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_5 = 4'hb == io_in_cnt ? 3'h4 : _GEN_70; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_6 = 4'hb == io_in_cnt ? 3'h7 : _GEN_82; // @[FFTDesigns.scala 3273:{17,17}]
endmodule
module PermutationsWithStreaming_6(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  input         io_in_en_5,
  input         io_in_en_6,
  input         io_in_en_7,
  input         io_in_en_8,
  input         io_in_en_9,
  input         io_in_en_10,
  input         io_in_en_11,
  input         io_in_en_12,
  input         io_in_en_13,
  input         io_in_en_14,
  input         io_in_en_15,
  input         io_in_en_16,
  input         io_in_en_17,
  input         io_in_en_18,
  input         io_in_en_19,
  input         io_in_en_20,
  input         io_in_en_21,
  input         io_in_en_22,
  input         io_in_en_23,
  input         io_in_en_24,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [4:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [4:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2641:26]
  wire [2:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [3:0] M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2642:27]
  wire [4:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2642:27]
  wire [4:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2642:27]
  wire [4:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2642:27]
  wire [4:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2642:27]
  wire [4:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2642:27]
  wire [4:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2642:27]
  wire [4:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2642:27]
  wire [4:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2643:27]
  wire [4:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2643:27]
  wire [4:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2643:27]
  wire [4:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2643:27]
  wire [4:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2643:27]
  wire [4:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2643:27]
  wire [4:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2643:27]
  wire [4:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2643:27]
  wire [4:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2643:27]
  wire [3:0] Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2644:29]
  wire [2:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2644:29]
  reg  offset_switch; // @[FFTDesigns.scala 2627:28]
  wire [5:0] lo_lo = {io_in_en_5,io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2628:19]
  wire [11:0] lo = {io_in_en_11,io_in_en_10,io_in_en_9,io_in_en_8,io_in_en_7,io_in_en_6,lo_lo}; // @[FFTDesigns.scala 2628:19]
  wire [5:0] hi_lo = {io_in_en_17,io_in_en_16,io_in_en_15,io_in_en_14,io_in_en_13,io_in_en_12}; // @[FFTDesigns.scala 2628:19]
  wire [24:0] _T = {io_in_en_24,io_in_en_23,io_in_en_22,io_in_en_21,io_in_en_20,io_in_en_19,io_in_en_18,hi_lo,lo}; // @[FFTDesigns.scala 2628:19]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2628:26]
  reg [3:0] cnt; // @[FFTDesigns.scala 2645:22]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2649:26]
  wire [3:0] _cnt_T_1 = cnt + 4'h1; // @[FFTDesigns.scala 2651:20]
  wire  _GEN_2 = cnt == 4'hb ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2647:32 2649:23 2652:23]
  wire [4:0] _T_6 = 4'hc * _offset_switch_T; // @[FFTDesigns.scala 2661:54]
  wire [4:0] _T_8 = M0_Config_ROM_io_out_0 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [4:0] _T_9 = 4'hc * offset_switch; // @[FFTDesigns.scala 2662:41]
  wire [4:0] _GEN_110 = {{1'd0}, cnt}; // @[FFTDesigns.scala 2662:31]
  wire [4:0] _T_11 = _GEN_110 + _T_9; // @[FFTDesigns.scala 2662:31]
  wire [4:0] _T_15 = _GEN_110 + _T_6; // @[FFTDesigns.scala 2664:31]
  wire [4:0] _T_18 = M1_Config_ROM_io_out_0 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [4:0] _T_22 = M0_Config_ROM_io_out_1 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [4:0] _T_32 = M1_Config_ROM_io_out_1 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [4:0] _T_36 = M0_Config_ROM_io_out_2 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [4:0] _T_46 = M1_Config_ROM_io_out_2 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [4:0] _T_50 = M0_Config_ROM_io_out_3 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [4:0] _T_60 = M1_Config_ROM_io_out_3 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [4:0] _T_64 = M0_Config_ROM_io_out_4 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [4:0] _T_74 = M1_Config_ROM_io_out_4 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [4:0] _T_78 = M0_Config_ROM_io_out_5 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [4:0] _T_88 = M1_Config_ROM_io_out_5 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [4:0] _T_92 = M0_Config_ROM_io_out_6 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [4:0] _T_102 = M1_Config_ROM_io_out_6 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [4:0] _T_106 = M0_Config_ROM_io_out_7 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [4:0] _T_116 = M1_Config_ROM_io_out_7 + _T_9; // @[FFTDesigns.scala 2665:44]
  RAM_Block_96 RAM_Block ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_1 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_2 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_3 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_4 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_5 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_6 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_7 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_8 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_9 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_10 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_11 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_12 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_13 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_14 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_15 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  PermutationModuleStreamed PermutationModuleStreamed ( // @[FFTDesigns.scala 2641:26]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im)
  );
  M0_Config_ROM_6 M0_Config_ROM ( // @[FFTDesigns.scala 2642:27]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7)
  );
  M1_Config_ROM_6 M1_Config_ROM ( // @[FFTDesigns.scala 2643:27]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7)
  );
  Streaming_Permute_Config_6 Streaming_Permute_Config ( // @[FFTDesigns.scala 2644:29]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6)
  );
  assign io_out_0_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_0_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = _T_1 ? _T_8 : 5'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_io_in_waddr = _T_1 ? _T_11 : 5'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_io_in_data_Re = io_in_0_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_in_data_Im = io_in_0_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = _T_1 ? _T_22 : 5'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_1_io_in_waddr = _T_1 ? _T_11 : 5'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_1_io_in_data_Re = io_in_1_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_in_data_Im = io_in_1_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = _T_1 ? _T_36 : 5'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_2_io_in_waddr = _T_1 ? _T_11 : 5'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_2_io_in_data_Re = io_in_2_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_in_data_Im = io_in_2_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = _T_1 ? _T_50 : 5'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_3_io_in_waddr = _T_1 ? _T_11 : 5'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_3_io_in_data_Re = io_in_3_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_in_data_Im = io_in_3_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = _T_1 ? _T_64 : 5'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_4_io_in_waddr = _T_1 ? _T_11 : 5'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_4_io_in_data_Re = io_in_4_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_in_data_Im = io_in_4_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = _T_1 ? _T_78 : 5'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_5_io_in_waddr = _T_1 ? _T_11 : 5'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_5_io_in_data_Re = io_in_5_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_in_data_Im = io_in_5_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = _T_1 ? _T_92 : 5'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_6_io_in_waddr = _T_1 ? _T_11 : 5'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_6_io_in_data_Re = io_in_6_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_in_data_Im = io_in_6_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = _T_1 ? _T_106 : 5'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_7_io_in_waddr = _T_1 ? _T_11 : 5'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_7_io_in_data_Re = io_in_7_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_in_data_Im = io_in_7_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = _T_1 ? _T_15 : 5'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_8_io_in_waddr = _T_1 ? _T_18 : 5'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_8_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_8_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = _T_1 ? _T_15 : 5'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_9_io_in_waddr = _T_1 ? _T_32 : 5'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_9_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_9_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = _T_1 ? _T_15 : 5'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_10_io_in_waddr = _T_1 ? _T_46 : 5'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_10_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_10_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = _T_1 ? _T_15 : 5'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_11_io_in_waddr = _T_1 ? _T_60 : 5'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_11_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_11_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = _T_1 ? _T_15 : 5'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_12_io_in_waddr = _T_1 ? _T_74 : 5'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_12_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_12_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = _T_1 ? _T_15 : 5'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_13_io_in_waddr = _T_1 ? _T_88 : 5'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_13_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_13_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = _T_1 ? _T_15 : 5'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_14_io_in_waddr = _T_1 ? _T_102 : 5'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_14_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_14_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = _T_1 ? _T_15 : 5'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_15_io_in_waddr = _T_1 ? _T_116 : 5'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_15_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_15_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign M0_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2694:22]
  assign M1_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2695:22]
  assign Streaming_Permute_Config_io_in_cnt = cnt; // @[FFTDesigns.scala 2696:24]
  always @(posedge clock) begin
    offset_switch <= _T_1 & _GEN_2; // @[FFTDesigns.scala 2646:30 2691:21]
    if (reset) begin // @[FFTDesigns.scala 2645:22]
      cnt <= 4'h0; // @[FFTDesigns.scala 2645:22]
    end else if (_T_1) begin // @[FFTDesigns.scala 2646:30]
      if (cnt == 4'hb) begin // @[FFTDesigns.scala 2647:32]
        cnt <= 4'h0; // @[FFTDesigns.scala 2648:13]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2651:13]
      end
    end else begin
      cnt <= 4'h0; // @[FFTDesigns.scala 2692:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_Block_112(
  input         clock,
  input  [3:0]  io_in_raddr,
  input  [3:0]  io_in_waddr,
  input  [31:0] io_in_data_Re,
  input  [31:0] io_in_data_Im,
  input         io_re,
  input         io_wr,
  input         io_en,
  output [31:0] io_out_data_Re,
  output [31:0] io_out_data_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_0_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_8_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_8_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_9_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_9_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_10_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_10_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_11_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_11_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_12_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_12_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_13_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_13_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_14_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_14_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_15_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_15_Im; // @[FFTDesigns.scala 3286:18]
  wire [31:0] _GEN_65 = 4'h1 == io_in_raddr ? mem_1_Im : mem_0_Im; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_66 = 4'h2 == io_in_raddr ? mem_2_Im : _GEN_65; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_67 = 4'h3 == io_in_raddr ? mem_3_Im : _GEN_66; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_68 = 4'h4 == io_in_raddr ? mem_4_Im : _GEN_67; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_69 = 4'h5 == io_in_raddr ? mem_5_Im : _GEN_68; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_70 = 4'h6 == io_in_raddr ? mem_6_Im : _GEN_69; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_71 = 4'h7 == io_in_raddr ? mem_7_Im : _GEN_70; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_72 = 4'h8 == io_in_raddr ? mem_8_Im : _GEN_71; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_73 = 4'h9 == io_in_raddr ? mem_9_Im : _GEN_72; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_74 = 4'ha == io_in_raddr ? mem_10_Im : _GEN_73; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_75 = 4'hb == io_in_raddr ? mem_11_Im : _GEN_74; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_76 = 4'hc == io_in_raddr ? mem_12_Im : _GEN_75; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_77 = 4'hd == io_in_raddr ? mem_13_Im : _GEN_76; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_78 = 4'he == io_in_raddr ? mem_14_Im : _GEN_77; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_79 = 4'hf == io_in_raddr ? mem_15_Im : _GEN_78; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_81 = 4'h1 == io_in_raddr ? mem_1_Re : mem_0_Re; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_82 = 4'h2 == io_in_raddr ? mem_2_Re : _GEN_81; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_83 = 4'h3 == io_in_raddr ? mem_3_Re : _GEN_82; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_84 = 4'h4 == io_in_raddr ? mem_4_Re : _GEN_83; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_85 = 4'h5 == io_in_raddr ? mem_5_Re : _GEN_84; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_86 = 4'h6 == io_in_raddr ? mem_6_Re : _GEN_85; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_87 = 4'h7 == io_in_raddr ? mem_7_Re : _GEN_86; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_88 = 4'h8 == io_in_raddr ? mem_8_Re : _GEN_87; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_89 = 4'h9 == io_in_raddr ? mem_9_Re : _GEN_88; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_90 = 4'ha == io_in_raddr ? mem_10_Re : _GEN_89; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_91 = 4'hb == io_in_raddr ? mem_11_Re : _GEN_90; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_92 = 4'hc == io_in_raddr ? mem_12_Re : _GEN_91; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_93 = 4'hd == io_in_raddr ? mem_13_Re : _GEN_92; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_94 = 4'he == io_in_raddr ? mem_14_Re : _GEN_93; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_95 = 4'hf == io_in_raddr ? mem_15_Re : _GEN_94; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_96 = io_re ? _GEN_79 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3295:24]
  wire [31:0] _GEN_97 = io_re ? _GEN_95 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3294:24]
  assign io_out_data_Re = io_en ? _GEN_97 : 32'h0; // @[FFTDesigns.scala 3287:16 3298:22]
  assign io_out_data_Im = io_en ? _GEN_96 : 32'h0; // @[FFTDesigns.scala 3287:16 3299:22]
  always @(posedge clock) begin
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h8 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_8_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h8 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_8_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h9 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_9_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h9 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_9_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'ha == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_10_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'ha == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_10_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hb == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_11_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hb == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_11_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hc == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_12_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hc == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_12_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hd == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_13_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hd == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_13_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'he == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_14_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'he == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_14_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hf == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_15_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hf == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_15_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_3_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_4_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_4_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_5_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_5_Im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_6_Re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_6_Im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_7_Re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_7_Im = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mem_8_Re = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mem_8_Im = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_9_Re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mem_9_Im = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mem_10_Re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mem_10_Im = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_11_Re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mem_11_Im = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  mem_12_Re = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  mem_12_Im = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  mem_13_Re = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mem_13_Im = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mem_14_Re = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mem_14_Im = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mem_15_Re = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mem_15_Im = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PermutationModuleStreamed_7(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [3:0]  io_in_config_0,
  input  [3:0]  io_in_config_1,
  input  [3:0]  io_in_config_2,
  input  [3:0]  io_in_config_3,
  input  [3:0]  io_in_config_4,
  input  [3:0]  io_in_config_5,
  input  [3:0]  io_in_config_6,
  input  [3:0]  io_in_config_7,
  input  [3:0]  io_in_config_8,
  input  [3:0]  io_in_config_9,
  input  [3:0]  io_in_config_10,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im
);
  wire  _T = io_in_config_0 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_1 = io_in_config_1 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_2 = io_in_config_2 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_3 = io_in_config_3 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_4 = io_in_config_4 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_5 = io_in_config_5 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_6 = io_in_config_6 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_7 = io_in_config_7 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_8 = io_in_config_8 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_9 = io_in_config_9 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_10 = io_in_config_10 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_12 = io_in_config_0 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_13 = io_in_config_1 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_14 = io_in_config_2 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_15 = io_in_config_3 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_16 = io_in_config_4 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_17 = io_in_config_5 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_18 = io_in_config_6 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_19 = io_in_config_7 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_20 = io_in_config_8 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_21 = io_in_config_9 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_22 = io_in_config_10 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_24 = io_in_config_0 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_25 = io_in_config_1 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_26 = io_in_config_2 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_27 = io_in_config_3 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_28 = io_in_config_4 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_29 = io_in_config_5 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_30 = io_in_config_6 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_31 = io_in_config_7 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_32 = io_in_config_8 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_33 = io_in_config_9 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_34 = io_in_config_10 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_36 = io_in_config_0 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_37 = io_in_config_1 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_38 = io_in_config_2 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_39 = io_in_config_3 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_40 = io_in_config_4 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_41 = io_in_config_5 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_42 = io_in_config_6 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_43 = io_in_config_7 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_44 = io_in_config_8 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_45 = io_in_config_9 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_46 = io_in_config_10 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_48 = io_in_config_0 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_49 = io_in_config_1 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_50 = io_in_config_2 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_51 = io_in_config_3 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_52 = io_in_config_4 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_53 = io_in_config_5 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_54 = io_in_config_6 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_55 = io_in_config_7 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_56 = io_in_config_8 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_57 = io_in_config_9 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_58 = io_in_config_10 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_60 = io_in_config_0 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_61 = io_in_config_1 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_62 = io_in_config_2 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_63 = io_in_config_3 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_64 = io_in_config_4 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_65 = io_in_config_5 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_66 = io_in_config_6 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_67 = io_in_config_7 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_68 = io_in_config_8 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_69 = io_in_config_9 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_70 = io_in_config_10 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_72 = io_in_config_0 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_73 = io_in_config_1 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_74 = io_in_config_2 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_75 = io_in_config_3 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_76 = io_in_config_4 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_77 = io_in_config_5 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_78 = io_in_config_6 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_79 = io_in_config_7 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_80 = io_in_config_8 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_81 = io_in_config_9 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_82 = io_in_config_10 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_84 = io_in_config_0 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_85 = io_in_config_1 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_86 = io_in_config_2 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_87 = io_in_config_3 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_88 = io_in_config_4 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_89 = io_in_config_5 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_90 = io_in_config_6 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_91 = io_in_config_7 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_92 = io_in_config_8 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_93 = io_in_config_9 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_94 = io_in_config_10 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_96 = io_in_config_0 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_97 = io_in_config_1 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_98 = io_in_config_2 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_99 = io_in_config_3 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_100 = io_in_config_4 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_101 = io_in_config_5 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_102 = io_in_config_6 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_103 = io_in_config_7 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_104 = io_in_config_8 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_105 = io_in_config_9 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_106 = io_in_config_10 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_108 = io_in_config_0 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_109 = io_in_config_1 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_110 = io_in_config_2 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_111 = io_in_config_3 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_112 = io_in_config_4 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_113 = io_in_config_5 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_114 = io_in_config_6 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_115 = io_in_config_7 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_116 = io_in_config_8 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_117 = io_in_config_9 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_118 = io_in_config_10 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_120 = io_in_config_0 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_121 = io_in_config_1 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_122 = io_in_config_2 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_123 = io_in_config_3 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_124 = io_in_config_4 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_125 = io_in_config_5 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_126 = io_in_config_6 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_127 = io_in_config_7 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_128 = io_in_config_8 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_129 = io_in_config_9 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_130 = io_in_config_10 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_132 = io_in_config_0 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_133 = io_in_config_1 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_134 = io_in_config_2 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_135 = io_in_config_3 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_136 = io_in_config_4 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_137 = io_in_config_5 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_138 = io_in_config_6 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_139 = io_in_config_7 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_140 = io_in_config_8 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_141 = io_in_config_9 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_142 = io_in_config_10 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire [3:0] _pms_pmx_T = _T_10 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_1 = _T_9 ? 4'h9 : _pms_pmx_T; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_2 = _T_8 ? 4'h8 : _pms_pmx_T_1; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_3 = _T_7 ? 4'h7 : _pms_pmx_T_2; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_4 = _T_6 ? 4'h6 : _pms_pmx_T_3; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_5 = _T_5 ? 4'h5 : _pms_pmx_T_4; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_6 = _T_4 ? 4'h4 : _pms_pmx_T_5; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_7 = _T_3 ? 4'h3 : _pms_pmx_T_6; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_8 = _T_2 ? 4'h2 : _pms_pmx_T_7; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_9 = _T_1 ? 4'h1 : _pms_pmx_T_8; // @[Mux.scala 47:70]
  wire [3:0] pms_0 = _T ? 4'h0 : _pms_pmx_T_9; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_10 = _T_22 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_11 = _T_21 ? 4'h9 : _pms_pmx_T_10; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_12 = _T_20 ? 4'h8 : _pms_pmx_T_11; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_13 = _T_19 ? 4'h7 : _pms_pmx_T_12; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_14 = _T_18 ? 4'h6 : _pms_pmx_T_13; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_15 = _T_17 ? 4'h5 : _pms_pmx_T_14; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_16 = _T_16 ? 4'h4 : _pms_pmx_T_15; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_17 = _T_15 ? 4'h3 : _pms_pmx_T_16; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_18 = _T_14 ? 4'h2 : _pms_pmx_T_17; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_19 = _T_13 ? 4'h1 : _pms_pmx_T_18; // @[Mux.scala 47:70]
  wire [3:0] pms_1 = _T_12 ? 4'h0 : _pms_pmx_T_19; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_20 = _T_34 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_21 = _T_33 ? 4'h9 : _pms_pmx_T_20; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_22 = _T_32 ? 4'h8 : _pms_pmx_T_21; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_23 = _T_31 ? 4'h7 : _pms_pmx_T_22; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_24 = _T_30 ? 4'h6 : _pms_pmx_T_23; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_25 = _T_29 ? 4'h5 : _pms_pmx_T_24; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_26 = _T_28 ? 4'h4 : _pms_pmx_T_25; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_27 = _T_27 ? 4'h3 : _pms_pmx_T_26; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_28 = _T_26 ? 4'h2 : _pms_pmx_T_27; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_29 = _T_25 ? 4'h1 : _pms_pmx_T_28; // @[Mux.scala 47:70]
  wire [3:0] pms_2 = _T_24 ? 4'h0 : _pms_pmx_T_29; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_30 = _T_46 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_31 = _T_45 ? 4'h9 : _pms_pmx_T_30; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_32 = _T_44 ? 4'h8 : _pms_pmx_T_31; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_33 = _T_43 ? 4'h7 : _pms_pmx_T_32; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_34 = _T_42 ? 4'h6 : _pms_pmx_T_33; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_35 = _T_41 ? 4'h5 : _pms_pmx_T_34; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_36 = _T_40 ? 4'h4 : _pms_pmx_T_35; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_37 = _T_39 ? 4'h3 : _pms_pmx_T_36; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_38 = _T_38 ? 4'h2 : _pms_pmx_T_37; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_39 = _T_37 ? 4'h1 : _pms_pmx_T_38; // @[Mux.scala 47:70]
  wire [3:0] pms_3 = _T_36 ? 4'h0 : _pms_pmx_T_39; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_40 = _T_58 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_41 = _T_57 ? 4'h9 : _pms_pmx_T_40; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_42 = _T_56 ? 4'h8 : _pms_pmx_T_41; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_43 = _T_55 ? 4'h7 : _pms_pmx_T_42; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_44 = _T_54 ? 4'h6 : _pms_pmx_T_43; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_45 = _T_53 ? 4'h5 : _pms_pmx_T_44; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_46 = _T_52 ? 4'h4 : _pms_pmx_T_45; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_47 = _T_51 ? 4'h3 : _pms_pmx_T_46; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_48 = _T_50 ? 4'h2 : _pms_pmx_T_47; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_49 = _T_49 ? 4'h1 : _pms_pmx_T_48; // @[Mux.scala 47:70]
  wire [3:0] pms_4 = _T_48 ? 4'h0 : _pms_pmx_T_49; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_50 = _T_70 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_51 = _T_69 ? 4'h9 : _pms_pmx_T_50; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_52 = _T_68 ? 4'h8 : _pms_pmx_T_51; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_53 = _T_67 ? 4'h7 : _pms_pmx_T_52; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_54 = _T_66 ? 4'h6 : _pms_pmx_T_53; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_55 = _T_65 ? 4'h5 : _pms_pmx_T_54; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_56 = _T_64 ? 4'h4 : _pms_pmx_T_55; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_57 = _T_63 ? 4'h3 : _pms_pmx_T_56; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_58 = _T_62 ? 4'h2 : _pms_pmx_T_57; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_59 = _T_61 ? 4'h1 : _pms_pmx_T_58; // @[Mux.scala 47:70]
  wire [3:0] pms_5 = _T_60 ? 4'h0 : _pms_pmx_T_59; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_60 = _T_82 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_61 = _T_81 ? 4'h9 : _pms_pmx_T_60; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_62 = _T_80 ? 4'h8 : _pms_pmx_T_61; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_63 = _T_79 ? 4'h7 : _pms_pmx_T_62; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_64 = _T_78 ? 4'h6 : _pms_pmx_T_63; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_65 = _T_77 ? 4'h5 : _pms_pmx_T_64; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_66 = _T_76 ? 4'h4 : _pms_pmx_T_65; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_67 = _T_75 ? 4'h3 : _pms_pmx_T_66; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_68 = _T_74 ? 4'h2 : _pms_pmx_T_67; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_69 = _T_73 ? 4'h1 : _pms_pmx_T_68; // @[Mux.scala 47:70]
  wire [3:0] pms_6 = _T_72 ? 4'h0 : _pms_pmx_T_69; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_70 = _T_94 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_71 = _T_93 ? 4'h9 : _pms_pmx_T_70; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_72 = _T_92 ? 4'h8 : _pms_pmx_T_71; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_73 = _T_91 ? 4'h7 : _pms_pmx_T_72; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_74 = _T_90 ? 4'h6 : _pms_pmx_T_73; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_75 = _T_89 ? 4'h5 : _pms_pmx_T_74; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_76 = _T_88 ? 4'h4 : _pms_pmx_T_75; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_77 = _T_87 ? 4'h3 : _pms_pmx_T_76; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_78 = _T_86 ? 4'h2 : _pms_pmx_T_77; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_79 = _T_85 ? 4'h1 : _pms_pmx_T_78; // @[Mux.scala 47:70]
  wire [3:0] pms_7 = _T_84 ? 4'h0 : _pms_pmx_T_79; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_80 = _T_106 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_81 = _T_105 ? 4'h9 : _pms_pmx_T_80; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_82 = _T_104 ? 4'h8 : _pms_pmx_T_81; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_83 = _T_103 ? 4'h7 : _pms_pmx_T_82; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_84 = _T_102 ? 4'h6 : _pms_pmx_T_83; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_85 = _T_101 ? 4'h5 : _pms_pmx_T_84; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_86 = _T_100 ? 4'h4 : _pms_pmx_T_85; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_87 = _T_99 ? 4'h3 : _pms_pmx_T_86; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_88 = _T_98 ? 4'h2 : _pms_pmx_T_87; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_89 = _T_97 ? 4'h1 : _pms_pmx_T_88; // @[Mux.scala 47:70]
  wire [3:0] pms_8 = _T_96 ? 4'h0 : _pms_pmx_T_89; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_90 = _T_118 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_91 = _T_117 ? 4'h9 : _pms_pmx_T_90; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_92 = _T_116 ? 4'h8 : _pms_pmx_T_91; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_93 = _T_115 ? 4'h7 : _pms_pmx_T_92; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_94 = _T_114 ? 4'h6 : _pms_pmx_T_93; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_95 = _T_113 ? 4'h5 : _pms_pmx_T_94; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_96 = _T_112 ? 4'h4 : _pms_pmx_T_95; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_97 = _T_111 ? 4'h3 : _pms_pmx_T_96; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_98 = _T_110 ? 4'h2 : _pms_pmx_T_97; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_99 = _T_109 ? 4'h1 : _pms_pmx_T_98; // @[Mux.scala 47:70]
  wire [3:0] pms_9 = _T_108 ? 4'h0 : _pms_pmx_T_99; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_100 = _T_130 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_101 = _T_129 ? 4'h9 : _pms_pmx_T_100; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_102 = _T_128 ? 4'h8 : _pms_pmx_T_101; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_103 = _T_127 ? 4'h7 : _pms_pmx_T_102; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_104 = _T_126 ? 4'h6 : _pms_pmx_T_103; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_105 = _T_125 ? 4'h5 : _pms_pmx_T_104; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_106 = _T_124 ? 4'h4 : _pms_pmx_T_105; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_107 = _T_123 ? 4'h3 : _pms_pmx_T_106; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_108 = _T_122 ? 4'h2 : _pms_pmx_T_107; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_109 = _T_121 ? 4'h1 : _pms_pmx_T_108; // @[Mux.scala 47:70]
  wire [3:0] pms_10 = _T_120 ? 4'h0 : _pms_pmx_T_109; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_110 = _T_142 ? 4'ha : 4'hb; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_111 = _T_141 ? 4'h9 : _pms_pmx_T_110; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_112 = _T_140 ? 4'h8 : _pms_pmx_T_111; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_113 = _T_139 ? 4'h7 : _pms_pmx_T_112; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_114 = _T_138 ? 4'h6 : _pms_pmx_T_113; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_115 = _T_137 ? 4'h5 : _pms_pmx_T_114; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_116 = _T_136 ? 4'h4 : _pms_pmx_T_115; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_117 = _T_135 ? 4'h3 : _pms_pmx_T_116; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_118 = _T_134 ? 4'h2 : _pms_pmx_T_117; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_119 = _T_133 ? 4'h1 : _pms_pmx_T_118; // @[Mux.scala 47:70]
  wire [3:0] pms_11 = _T_132 ? 4'h0 : _pms_pmx_T_119; // @[Mux.scala 47:70]
  wire [31:0] _GEN_1 = 4'h1 == pms_0 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_2 = 4'h2 == pms_0 ? io_in_2_Im : _GEN_1; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_3 = 4'h3 == pms_0 ? io_in_3_Im : _GEN_2; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_4 = 4'h4 == pms_0 ? io_in_4_Im : _GEN_3; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_5 = 4'h5 == pms_0 ? io_in_5_Im : _GEN_4; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_6 = 4'h6 == pms_0 ? io_in_6_Im : _GEN_5; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_7 = 4'h7 == pms_0 ? io_in_7_Im : _GEN_6; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_8 = 4'h8 == pms_0 ? io_in_8_Im : _GEN_7; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_9 = 4'h9 == pms_0 ? io_in_9_Im : _GEN_8; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_10 = 4'ha == pms_0 ? io_in_10_Im : _GEN_9; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_13 = 4'h1 == pms_0 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_14 = 4'h2 == pms_0 ? io_in_2_Re : _GEN_13; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_15 = 4'h3 == pms_0 ? io_in_3_Re : _GEN_14; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_16 = 4'h4 == pms_0 ? io_in_4_Re : _GEN_15; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_17 = 4'h5 == pms_0 ? io_in_5_Re : _GEN_16; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_18 = 4'h6 == pms_0 ? io_in_6_Re : _GEN_17; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_19 = 4'h7 == pms_0 ? io_in_7_Re : _GEN_18; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_20 = 4'h8 == pms_0 ? io_in_8_Re : _GEN_19; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_21 = 4'h9 == pms_0 ? io_in_9_Re : _GEN_20; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_22 = 4'ha == pms_0 ? io_in_10_Re : _GEN_21; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_25 = 4'h1 == pms_1 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_26 = 4'h2 == pms_1 ? io_in_2_Im : _GEN_25; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_27 = 4'h3 == pms_1 ? io_in_3_Im : _GEN_26; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_28 = 4'h4 == pms_1 ? io_in_4_Im : _GEN_27; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_29 = 4'h5 == pms_1 ? io_in_5_Im : _GEN_28; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_30 = 4'h6 == pms_1 ? io_in_6_Im : _GEN_29; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_31 = 4'h7 == pms_1 ? io_in_7_Im : _GEN_30; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_32 = 4'h8 == pms_1 ? io_in_8_Im : _GEN_31; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_33 = 4'h9 == pms_1 ? io_in_9_Im : _GEN_32; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_34 = 4'ha == pms_1 ? io_in_10_Im : _GEN_33; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_37 = 4'h1 == pms_1 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_38 = 4'h2 == pms_1 ? io_in_2_Re : _GEN_37; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_39 = 4'h3 == pms_1 ? io_in_3_Re : _GEN_38; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_40 = 4'h4 == pms_1 ? io_in_4_Re : _GEN_39; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_41 = 4'h5 == pms_1 ? io_in_5_Re : _GEN_40; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_42 = 4'h6 == pms_1 ? io_in_6_Re : _GEN_41; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_43 = 4'h7 == pms_1 ? io_in_7_Re : _GEN_42; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_44 = 4'h8 == pms_1 ? io_in_8_Re : _GEN_43; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_45 = 4'h9 == pms_1 ? io_in_9_Re : _GEN_44; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_46 = 4'ha == pms_1 ? io_in_10_Re : _GEN_45; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_49 = 4'h1 == pms_2 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_50 = 4'h2 == pms_2 ? io_in_2_Im : _GEN_49; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_51 = 4'h3 == pms_2 ? io_in_3_Im : _GEN_50; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_52 = 4'h4 == pms_2 ? io_in_4_Im : _GEN_51; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_53 = 4'h5 == pms_2 ? io_in_5_Im : _GEN_52; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_54 = 4'h6 == pms_2 ? io_in_6_Im : _GEN_53; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_55 = 4'h7 == pms_2 ? io_in_7_Im : _GEN_54; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_56 = 4'h8 == pms_2 ? io_in_8_Im : _GEN_55; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_57 = 4'h9 == pms_2 ? io_in_9_Im : _GEN_56; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_58 = 4'ha == pms_2 ? io_in_10_Im : _GEN_57; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_61 = 4'h1 == pms_2 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_62 = 4'h2 == pms_2 ? io_in_2_Re : _GEN_61; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_63 = 4'h3 == pms_2 ? io_in_3_Re : _GEN_62; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_64 = 4'h4 == pms_2 ? io_in_4_Re : _GEN_63; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_65 = 4'h5 == pms_2 ? io_in_5_Re : _GEN_64; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_66 = 4'h6 == pms_2 ? io_in_6_Re : _GEN_65; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_67 = 4'h7 == pms_2 ? io_in_7_Re : _GEN_66; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_68 = 4'h8 == pms_2 ? io_in_8_Re : _GEN_67; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_69 = 4'h9 == pms_2 ? io_in_9_Re : _GEN_68; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_70 = 4'ha == pms_2 ? io_in_10_Re : _GEN_69; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_73 = 4'h1 == pms_3 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_74 = 4'h2 == pms_3 ? io_in_2_Im : _GEN_73; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_75 = 4'h3 == pms_3 ? io_in_3_Im : _GEN_74; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_76 = 4'h4 == pms_3 ? io_in_4_Im : _GEN_75; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_77 = 4'h5 == pms_3 ? io_in_5_Im : _GEN_76; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_78 = 4'h6 == pms_3 ? io_in_6_Im : _GEN_77; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_79 = 4'h7 == pms_3 ? io_in_7_Im : _GEN_78; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_80 = 4'h8 == pms_3 ? io_in_8_Im : _GEN_79; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_81 = 4'h9 == pms_3 ? io_in_9_Im : _GEN_80; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_82 = 4'ha == pms_3 ? io_in_10_Im : _GEN_81; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_85 = 4'h1 == pms_3 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_86 = 4'h2 == pms_3 ? io_in_2_Re : _GEN_85; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_87 = 4'h3 == pms_3 ? io_in_3_Re : _GEN_86; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_88 = 4'h4 == pms_3 ? io_in_4_Re : _GEN_87; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_89 = 4'h5 == pms_3 ? io_in_5_Re : _GEN_88; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_90 = 4'h6 == pms_3 ? io_in_6_Re : _GEN_89; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_91 = 4'h7 == pms_3 ? io_in_7_Re : _GEN_90; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_92 = 4'h8 == pms_3 ? io_in_8_Re : _GEN_91; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_93 = 4'h9 == pms_3 ? io_in_9_Re : _GEN_92; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_94 = 4'ha == pms_3 ? io_in_10_Re : _GEN_93; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_97 = 4'h1 == pms_4 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_98 = 4'h2 == pms_4 ? io_in_2_Im : _GEN_97; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_99 = 4'h3 == pms_4 ? io_in_3_Im : _GEN_98; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_100 = 4'h4 == pms_4 ? io_in_4_Im : _GEN_99; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_101 = 4'h5 == pms_4 ? io_in_5_Im : _GEN_100; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_102 = 4'h6 == pms_4 ? io_in_6_Im : _GEN_101; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_103 = 4'h7 == pms_4 ? io_in_7_Im : _GEN_102; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_104 = 4'h8 == pms_4 ? io_in_8_Im : _GEN_103; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_105 = 4'h9 == pms_4 ? io_in_9_Im : _GEN_104; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_106 = 4'ha == pms_4 ? io_in_10_Im : _GEN_105; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_109 = 4'h1 == pms_4 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_110 = 4'h2 == pms_4 ? io_in_2_Re : _GEN_109; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_111 = 4'h3 == pms_4 ? io_in_3_Re : _GEN_110; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_112 = 4'h4 == pms_4 ? io_in_4_Re : _GEN_111; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_113 = 4'h5 == pms_4 ? io_in_5_Re : _GEN_112; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_114 = 4'h6 == pms_4 ? io_in_6_Re : _GEN_113; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_115 = 4'h7 == pms_4 ? io_in_7_Re : _GEN_114; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_116 = 4'h8 == pms_4 ? io_in_8_Re : _GEN_115; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_117 = 4'h9 == pms_4 ? io_in_9_Re : _GEN_116; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_118 = 4'ha == pms_4 ? io_in_10_Re : _GEN_117; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_121 = 4'h1 == pms_5 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_122 = 4'h2 == pms_5 ? io_in_2_Im : _GEN_121; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_123 = 4'h3 == pms_5 ? io_in_3_Im : _GEN_122; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_124 = 4'h4 == pms_5 ? io_in_4_Im : _GEN_123; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_125 = 4'h5 == pms_5 ? io_in_5_Im : _GEN_124; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_126 = 4'h6 == pms_5 ? io_in_6_Im : _GEN_125; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_127 = 4'h7 == pms_5 ? io_in_7_Im : _GEN_126; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_128 = 4'h8 == pms_5 ? io_in_8_Im : _GEN_127; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_129 = 4'h9 == pms_5 ? io_in_9_Im : _GEN_128; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_130 = 4'ha == pms_5 ? io_in_10_Im : _GEN_129; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_133 = 4'h1 == pms_5 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_134 = 4'h2 == pms_5 ? io_in_2_Re : _GEN_133; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_135 = 4'h3 == pms_5 ? io_in_3_Re : _GEN_134; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_136 = 4'h4 == pms_5 ? io_in_4_Re : _GEN_135; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_137 = 4'h5 == pms_5 ? io_in_5_Re : _GEN_136; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_138 = 4'h6 == pms_5 ? io_in_6_Re : _GEN_137; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_139 = 4'h7 == pms_5 ? io_in_7_Re : _GEN_138; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_140 = 4'h8 == pms_5 ? io_in_8_Re : _GEN_139; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_141 = 4'h9 == pms_5 ? io_in_9_Re : _GEN_140; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_142 = 4'ha == pms_5 ? io_in_10_Re : _GEN_141; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_145 = 4'h1 == pms_6 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_146 = 4'h2 == pms_6 ? io_in_2_Im : _GEN_145; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_147 = 4'h3 == pms_6 ? io_in_3_Im : _GEN_146; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_148 = 4'h4 == pms_6 ? io_in_4_Im : _GEN_147; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_149 = 4'h5 == pms_6 ? io_in_5_Im : _GEN_148; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_150 = 4'h6 == pms_6 ? io_in_6_Im : _GEN_149; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_151 = 4'h7 == pms_6 ? io_in_7_Im : _GEN_150; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_152 = 4'h8 == pms_6 ? io_in_8_Im : _GEN_151; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_153 = 4'h9 == pms_6 ? io_in_9_Im : _GEN_152; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_154 = 4'ha == pms_6 ? io_in_10_Im : _GEN_153; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_157 = 4'h1 == pms_6 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_158 = 4'h2 == pms_6 ? io_in_2_Re : _GEN_157; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_159 = 4'h3 == pms_6 ? io_in_3_Re : _GEN_158; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_160 = 4'h4 == pms_6 ? io_in_4_Re : _GEN_159; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_161 = 4'h5 == pms_6 ? io_in_5_Re : _GEN_160; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_162 = 4'h6 == pms_6 ? io_in_6_Re : _GEN_161; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_163 = 4'h7 == pms_6 ? io_in_7_Re : _GEN_162; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_164 = 4'h8 == pms_6 ? io_in_8_Re : _GEN_163; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_165 = 4'h9 == pms_6 ? io_in_9_Re : _GEN_164; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_166 = 4'ha == pms_6 ? io_in_10_Re : _GEN_165; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_169 = 4'h1 == pms_7 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_170 = 4'h2 == pms_7 ? io_in_2_Im : _GEN_169; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_171 = 4'h3 == pms_7 ? io_in_3_Im : _GEN_170; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_172 = 4'h4 == pms_7 ? io_in_4_Im : _GEN_171; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_173 = 4'h5 == pms_7 ? io_in_5_Im : _GEN_172; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_174 = 4'h6 == pms_7 ? io_in_6_Im : _GEN_173; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_175 = 4'h7 == pms_7 ? io_in_7_Im : _GEN_174; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_176 = 4'h8 == pms_7 ? io_in_8_Im : _GEN_175; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_177 = 4'h9 == pms_7 ? io_in_9_Im : _GEN_176; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_178 = 4'ha == pms_7 ? io_in_10_Im : _GEN_177; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_181 = 4'h1 == pms_7 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_182 = 4'h2 == pms_7 ? io_in_2_Re : _GEN_181; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_183 = 4'h3 == pms_7 ? io_in_3_Re : _GEN_182; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_184 = 4'h4 == pms_7 ? io_in_4_Re : _GEN_183; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_185 = 4'h5 == pms_7 ? io_in_5_Re : _GEN_184; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_186 = 4'h6 == pms_7 ? io_in_6_Re : _GEN_185; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_187 = 4'h7 == pms_7 ? io_in_7_Re : _GEN_186; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_188 = 4'h8 == pms_7 ? io_in_8_Re : _GEN_187; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_189 = 4'h9 == pms_7 ? io_in_9_Re : _GEN_188; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_190 = 4'ha == pms_7 ? io_in_10_Re : _GEN_189; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_193 = 4'h1 == pms_8 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_194 = 4'h2 == pms_8 ? io_in_2_Im : _GEN_193; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_195 = 4'h3 == pms_8 ? io_in_3_Im : _GEN_194; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_196 = 4'h4 == pms_8 ? io_in_4_Im : _GEN_195; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_197 = 4'h5 == pms_8 ? io_in_5_Im : _GEN_196; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_198 = 4'h6 == pms_8 ? io_in_6_Im : _GEN_197; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_199 = 4'h7 == pms_8 ? io_in_7_Im : _GEN_198; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_200 = 4'h8 == pms_8 ? io_in_8_Im : _GEN_199; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_201 = 4'h9 == pms_8 ? io_in_9_Im : _GEN_200; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_202 = 4'ha == pms_8 ? io_in_10_Im : _GEN_201; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_205 = 4'h1 == pms_8 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_206 = 4'h2 == pms_8 ? io_in_2_Re : _GEN_205; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_207 = 4'h3 == pms_8 ? io_in_3_Re : _GEN_206; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_208 = 4'h4 == pms_8 ? io_in_4_Re : _GEN_207; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_209 = 4'h5 == pms_8 ? io_in_5_Re : _GEN_208; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_210 = 4'h6 == pms_8 ? io_in_6_Re : _GEN_209; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_211 = 4'h7 == pms_8 ? io_in_7_Re : _GEN_210; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_212 = 4'h8 == pms_8 ? io_in_8_Re : _GEN_211; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_213 = 4'h9 == pms_8 ? io_in_9_Re : _GEN_212; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_214 = 4'ha == pms_8 ? io_in_10_Re : _GEN_213; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_217 = 4'h1 == pms_9 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_218 = 4'h2 == pms_9 ? io_in_2_Im : _GEN_217; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_219 = 4'h3 == pms_9 ? io_in_3_Im : _GEN_218; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_220 = 4'h4 == pms_9 ? io_in_4_Im : _GEN_219; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_221 = 4'h5 == pms_9 ? io_in_5_Im : _GEN_220; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_222 = 4'h6 == pms_9 ? io_in_6_Im : _GEN_221; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_223 = 4'h7 == pms_9 ? io_in_7_Im : _GEN_222; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_224 = 4'h8 == pms_9 ? io_in_8_Im : _GEN_223; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_225 = 4'h9 == pms_9 ? io_in_9_Im : _GEN_224; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_226 = 4'ha == pms_9 ? io_in_10_Im : _GEN_225; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_229 = 4'h1 == pms_9 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_230 = 4'h2 == pms_9 ? io_in_2_Re : _GEN_229; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_231 = 4'h3 == pms_9 ? io_in_3_Re : _GEN_230; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_232 = 4'h4 == pms_9 ? io_in_4_Re : _GEN_231; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_233 = 4'h5 == pms_9 ? io_in_5_Re : _GEN_232; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_234 = 4'h6 == pms_9 ? io_in_6_Re : _GEN_233; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_235 = 4'h7 == pms_9 ? io_in_7_Re : _GEN_234; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_236 = 4'h8 == pms_9 ? io_in_8_Re : _GEN_235; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_237 = 4'h9 == pms_9 ? io_in_9_Re : _GEN_236; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_238 = 4'ha == pms_9 ? io_in_10_Re : _GEN_237; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_241 = 4'h1 == pms_10 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_242 = 4'h2 == pms_10 ? io_in_2_Im : _GEN_241; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_243 = 4'h3 == pms_10 ? io_in_3_Im : _GEN_242; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_244 = 4'h4 == pms_10 ? io_in_4_Im : _GEN_243; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_245 = 4'h5 == pms_10 ? io_in_5_Im : _GEN_244; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_246 = 4'h6 == pms_10 ? io_in_6_Im : _GEN_245; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_247 = 4'h7 == pms_10 ? io_in_7_Im : _GEN_246; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_248 = 4'h8 == pms_10 ? io_in_8_Im : _GEN_247; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_249 = 4'h9 == pms_10 ? io_in_9_Im : _GEN_248; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_250 = 4'ha == pms_10 ? io_in_10_Im : _GEN_249; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_253 = 4'h1 == pms_10 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_254 = 4'h2 == pms_10 ? io_in_2_Re : _GEN_253; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_255 = 4'h3 == pms_10 ? io_in_3_Re : _GEN_254; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_256 = 4'h4 == pms_10 ? io_in_4_Re : _GEN_255; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_257 = 4'h5 == pms_10 ? io_in_5_Re : _GEN_256; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_258 = 4'h6 == pms_10 ? io_in_6_Re : _GEN_257; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_259 = 4'h7 == pms_10 ? io_in_7_Re : _GEN_258; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_260 = 4'h8 == pms_10 ? io_in_8_Re : _GEN_259; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_261 = 4'h9 == pms_10 ? io_in_9_Re : _GEN_260; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_262 = 4'ha == pms_10 ? io_in_10_Re : _GEN_261; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_265 = 4'h1 == pms_11 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_266 = 4'h2 == pms_11 ? io_in_2_Im : _GEN_265; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_267 = 4'h3 == pms_11 ? io_in_3_Im : _GEN_266; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_268 = 4'h4 == pms_11 ? io_in_4_Im : _GEN_267; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_269 = 4'h5 == pms_11 ? io_in_5_Im : _GEN_268; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_270 = 4'h6 == pms_11 ? io_in_6_Im : _GEN_269; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_271 = 4'h7 == pms_11 ? io_in_7_Im : _GEN_270; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_272 = 4'h8 == pms_11 ? io_in_8_Im : _GEN_271; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_273 = 4'h9 == pms_11 ? io_in_9_Im : _GEN_272; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_274 = 4'ha == pms_11 ? io_in_10_Im : _GEN_273; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_277 = 4'h1 == pms_11 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_278 = 4'h2 == pms_11 ? io_in_2_Re : _GEN_277; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_279 = 4'h3 == pms_11 ? io_in_3_Re : _GEN_278; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_280 = 4'h4 == pms_11 ? io_in_4_Re : _GEN_279; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_281 = 4'h5 == pms_11 ? io_in_5_Re : _GEN_280; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_282 = 4'h6 == pms_11 ? io_in_6_Re : _GEN_281; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_283 = 4'h7 == pms_11 ? io_in_7_Re : _GEN_282; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_284 = 4'h8 == pms_11 ? io_in_8_Re : _GEN_283; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_285 = 4'h9 == pms_11 ? io_in_9_Re : _GEN_284; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_286 = 4'ha == pms_11 ? io_in_10_Re : _GEN_285; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_0_Re = 4'hb == pms_0 ? io_in_11_Re : _GEN_22; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_0_Im = 4'hb == pms_0 ? io_in_11_Im : _GEN_10; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_1_Re = 4'hb == pms_1 ? io_in_11_Re : _GEN_46; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_1_Im = 4'hb == pms_1 ? io_in_11_Im : _GEN_34; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_2_Re = 4'hb == pms_2 ? io_in_11_Re : _GEN_70; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_2_Im = 4'hb == pms_2 ? io_in_11_Im : _GEN_58; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_3_Re = 4'hb == pms_3 ? io_in_11_Re : _GEN_94; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_3_Im = 4'hb == pms_3 ? io_in_11_Im : _GEN_82; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_4_Re = 4'hb == pms_4 ? io_in_11_Re : _GEN_118; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_4_Im = 4'hb == pms_4 ? io_in_11_Im : _GEN_106; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_5_Re = 4'hb == pms_5 ? io_in_11_Re : _GEN_142; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_5_Im = 4'hb == pms_5 ? io_in_11_Im : _GEN_130; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_6_Re = 4'hb == pms_6 ? io_in_11_Re : _GEN_166; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_6_Im = 4'hb == pms_6 ? io_in_11_Im : _GEN_154; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_7_Re = 4'hb == pms_7 ? io_in_11_Re : _GEN_190; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_7_Im = 4'hb == pms_7 ? io_in_11_Im : _GEN_178; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_8_Re = 4'hb == pms_8 ? io_in_11_Re : _GEN_214; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_8_Im = 4'hb == pms_8 ? io_in_11_Im : _GEN_202; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_9_Re = 4'hb == pms_9 ? io_in_11_Re : _GEN_238; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_9_Im = 4'hb == pms_9 ? io_in_11_Im : _GEN_226; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_10_Re = 4'hb == pms_10 ? io_in_11_Re : _GEN_262; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_10_Im = 4'hb == pms_10 ? io_in_11_Im : _GEN_250; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_11_Re = 4'hb == pms_11 ? io_in_11_Re : _GEN_286; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_11_Im = 4'hb == pms_11 ? io_in_11_Im : _GEN_274; // @[FFTDesigns.scala 3203:{17,17}]
endmodule
module M0_Config_ROM_7(
  input  [2:0] io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11
);
  wire [3:0] _GEN_1 = 3'h1 == io_in_cnt ? 4'h1 : 4'h0; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_2 = 3'h2 == io_in_cnt ? 4'h2 : _GEN_1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_3 = 3'h3 == io_in_cnt ? 4'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_4 = 3'h4 == io_in_cnt ? 4'h4 : _GEN_3; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_5 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_4; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_6 = 3'h6 == io_in_cnt ? 4'h6 : _GEN_5; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_33 = 3'h1 == io_in_cnt ? 4'h4 : 4'h3; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_34 = 3'h2 == io_in_cnt ? 4'h5 : _GEN_33; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_35 = 3'h3 == io_in_cnt ? 4'h6 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_36 = 3'h4 == io_in_cnt ? 4'h7 : _GEN_35; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_37 = 3'h5 == io_in_cnt ? 4'h0 : _GEN_36; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_38 = 3'h6 == io_in_cnt ? 4'h1 : _GEN_37; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_65 = 3'h1 == io_in_cnt ? 4'h6 : 4'h5; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_66 = 3'h2 == io_in_cnt ? 4'h2 : _GEN_65; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_67 = 3'h3 == io_in_cnt ? 4'h0 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_68 = 3'h4 == io_in_cnt ? 4'h1 : _GEN_67; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_69 = 3'h5 == io_in_cnt ? 4'h7 : _GEN_68; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_70 = 3'h6 == io_in_cnt ? 4'h3 : _GEN_69; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_0 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_1 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_2 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_3 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_6; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_4 = 3'h7 == io_in_cnt ? 4'h2 : _GEN_38; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_5 = 3'h7 == io_in_cnt ? 4'h2 : _GEN_38; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_6 = 3'h7 == io_in_cnt ? 4'h2 : _GEN_38; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_7 = 3'h7 == io_in_cnt ? 4'h2 : _GEN_38; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_8 = 3'h7 == io_in_cnt ? 4'h4 : _GEN_70; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_9 = 3'h7 == io_in_cnt ? 4'h4 : _GEN_70; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_10 = 3'h7 == io_in_cnt ? 4'h4 : _GEN_70; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_11 = 3'h7 == io_in_cnt ? 4'h4 : _GEN_70; // @[FFTDesigns.scala 3227:{17,17}]
endmodule
module M1_Config_ROM_7(
  input  [2:0] io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11
);
  wire [3:0] _GEN_1 = 3'h1 == io_in_cnt ? 4'h3 : 4'h0; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_2 = 3'h2 == io_in_cnt ? 4'h6 : _GEN_1; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_3 = 3'h3 == io_in_cnt ? 4'h2 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_4 = 3'h4 == io_in_cnt ? 4'h5 : _GEN_3; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_5 = 3'h5 == io_in_cnt ? 4'h1 : _GEN_4; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_6 = 3'h6 == io_in_cnt ? 4'h4 : _GEN_5; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_9 = 3'h1 == io_in_cnt ? 4'h5 : 4'h2; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_10 = 3'h2 == io_in_cnt ? 4'h0 : _GEN_9; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_11 = 3'h3 == io_in_cnt ? 4'h1 : _GEN_10; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_12 = 3'h4 == io_in_cnt ? 4'h4 : _GEN_11; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_13 = 3'h5 == io_in_cnt ? 4'h7 : _GEN_12; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_14 = 3'h6 == io_in_cnt ? 4'h3 : _GEN_13; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_17 = 3'h1 == io_in_cnt ? 4'h4 : 4'h1; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_18 = 3'h2 == io_in_cnt ? 4'h0 : _GEN_17; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_19 = 3'h3 == io_in_cnt ? 4'h3 : _GEN_18; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_20 = 3'h4 == io_in_cnt ? 4'h6 : _GEN_19; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_21 = 3'h5 == io_in_cnt ? 4'h7 : _GEN_20; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_22 = 3'h6 == io_in_cnt ? 4'h2 : _GEN_21; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_0 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_6; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_1 = 3'h7 == io_in_cnt ? 4'h6 : _GEN_14; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_2 = 3'h7 == io_in_cnt ? 4'h5 : _GEN_22; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_3 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_6; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_4 = 3'h7 == io_in_cnt ? 4'h6 : _GEN_14; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_5 = 3'h7 == io_in_cnt ? 4'h5 : _GEN_22; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_6 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_6; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_7 = 3'h7 == io_in_cnt ? 4'h6 : _GEN_14; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_8 = 3'h7 == io_in_cnt ? 4'h5 : _GEN_22; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_9 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_6; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_10 = 3'h7 == io_in_cnt ? 4'h6 : _GEN_14; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_11 = 3'h7 == io_in_cnt ? 4'h5 : _GEN_22; // @[FFTDesigns.scala 3250:{17,17}]
endmodule
module Streaming_Permute_Config_7(
  input  [2:0] io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10
);
  wire [3:0] _GEN_3 = 3'h3 == io_in_cnt ? 4'h1 : 4'h0; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_4 = 3'h4 == io_in_cnt ? 4'h1 : _GEN_3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_5 = 3'h5 == io_in_cnt ? 4'h1 : _GEN_4; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_6 = 3'h6 == io_in_cnt ? 4'h2 : _GEN_5; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_11 = 3'h3 == io_in_cnt ? 4'h4 : 4'h3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_12 = 3'h4 == io_in_cnt ? 4'h4 : _GEN_11; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_13 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_12; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_14 = 3'h6 == io_in_cnt ? 4'h5 : _GEN_13; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_19 = 3'h3 == io_in_cnt ? 4'h7 : 4'h6; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_20 = 3'h4 == io_in_cnt ? 4'h7 : _GEN_19; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_21 = 3'h5 == io_in_cnt ? 4'h7 : _GEN_20; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_22 = 3'h6 == io_in_cnt ? 4'h8 : _GEN_21; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_27 = 3'h3 == io_in_cnt ? 4'ha : 4'h9; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_28 = 3'h4 == io_in_cnt ? 4'ha : _GEN_27; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_29 = 3'h5 == io_in_cnt ? 4'ha : _GEN_28; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_30 = 3'h6 == io_in_cnt ? 4'hb : _GEN_29; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_34 = 3'h2 == io_in_cnt ? 4'h2 : 4'h1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_35 = 3'h3 == io_in_cnt ? 4'h2 : _GEN_34; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_36 = 3'h4 == io_in_cnt ? 4'h2 : _GEN_35; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_37 = 3'h5 == io_in_cnt ? 4'h0 : _GEN_36; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_38 = 3'h6 == io_in_cnt ? 4'h0 : _GEN_37; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_42 = 3'h2 == io_in_cnt ? 4'h5 : 4'h4; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_43 = 3'h3 == io_in_cnt ? 4'h5 : _GEN_42; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_44 = 3'h4 == io_in_cnt ? 4'h5 : _GEN_43; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_45 = 3'h5 == io_in_cnt ? 4'h3 : _GEN_44; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_46 = 3'h6 == io_in_cnt ? 4'h3 : _GEN_45; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_50 = 3'h2 == io_in_cnt ? 4'h8 : 4'h7; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_51 = 3'h3 == io_in_cnt ? 4'h8 : _GEN_50; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_52 = 3'h4 == io_in_cnt ? 4'h8 : _GEN_51; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_53 = 3'h5 == io_in_cnt ? 4'h6 : _GEN_52; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_54 = 3'h6 == io_in_cnt ? 4'h6 : _GEN_53; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_58 = 3'h2 == io_in_cnt ? 4'hb : 4'ha; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_59 = 3'h3 == io_in_cnt ? 4'hb : _GEN_58; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_60 = 3'h4 == io_in_cnt ? 4'hb : _GEN_59; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_61 = 3'h5 == io_in_cnt ? 4'h9 : _GEN_60; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_62 = 3'h6 == io_in_cnt ? 4'h9 : _GEN_61; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_66 = 3'h2 == io_in_cnt ? 4'h1 : 4'h2; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_67 = 3'h3 == io_in_cnt ? 4'h0 : _GEN_66; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_68 = 3'h4 == io_in_cnt ? 4'h0 : _GEN_67; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_69 = 3'h5 == io_in_cnt ? 4'h2 : _GEN_68; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_70 = 3'h6 == io_in_cnt ? 4'h1 : _GEN_69; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_74 = 3'h2 == io_in_cnt ? 4'h4 : 4'h5; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_75 = 3'h3 == io_in_cnt ? 4'h3 : _GEN_74; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_76 = 3'h4 == io_in_cnt ? 4'h3 : _GEN_75; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_77 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_76; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_78 = 3'h6 == io_in_cnt ? 4'h4 : _GEN_77; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_82 = 3'h2 == io_in_cnt ? 4'h7 : 4'h8; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_83 = 3'h3 == io_in_cnt ? 4'h6 : _GEN_82; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_84 = 3'h4 == io_in_cnt ? 4'h6 : _GEN_83; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_85 = 3'h5 == io_in_cnt ? 4'h8 : _GEN_84; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_86 = 3'h6 == io_in_cnt ? 4'h7 : _GEN_85; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_0 = 3'h7 == io_in_cnt ? 4'h2 : _GEN_6; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_1 = 3'h7 == io_in_cnt ? 4'h5 : _GEN_14; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_2 = 3'h7 == io_in_cnt ? 4'h8 : _GEN_22; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_3 = 3'h7 == io_in_cnt ? 4'hb : _GEN_30; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_4 = 3'h7 == io_in_cnt ? 4'h0 : _GEN_38; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_5 = 3'h7 == io_in_cnt ? 4'h3 : _GEN_46; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_6 = 3'h7 == io_in_cnt ? 4'h6 : _GEN_54; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_7 = 3'h7 == io_in_cnt ? 4'h9 : _GEN_62; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_8 = 3'h7 == io_in_cnt ? 4'h1 : _GEN_70; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_9 = 3'h7 == io_in_cnt ? 4'h4 : _GEN_78; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_10 = 3'h7 == io_in_cnt ? 4'h7 : _GEN_86; // @[FFTDesigns.scala 3273:{17,17}]
endmodule
module PermutationsWithStreaming_mr(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  input         io_in_en_5,
  input         io_in_en_6,
  input         io_in_en_7,
  input         io_in_en_8,
  input         io_in_en_9,
  input         io_in_en_10,
  input         io_in_en_11,
  input         io_in_en_12,
  input         io_in_en_13,
  input         io_in_en_14,
  input         io_in_en_15,
  input         io_in_en_16,
  input         io_in_en_17,
  input         io_in_en_18,
  input         io_in_en_19,
  input         io_in_en_20,
  input         io_in_en_21,
  input         io_in_en_22,
  input         io_in_en_23,
  input         io_in_en_24,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [3:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_16_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_16_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_16_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_16_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_16_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_16_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_16_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_16_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_17_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_17_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_17_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_17_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_17_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_17_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_17_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_17_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_18_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_18_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_18_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_18_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_18_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_18_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_18_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_18_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_19_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_19_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_19_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_19_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_19_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_19_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_19_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_19_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_20_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_20_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_20_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_20_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_20_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_20_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_20_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_20_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_21_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_21_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_21_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_21_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_21_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_21_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_21_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_21_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_22_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_22_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_22_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_22_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_22_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_22_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_22_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_22_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_23_clock; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_23_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [3:0] RAM_Block_23_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_23_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_23_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_23_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_23_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_23_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_8_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_8_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_9_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_9_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_10_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_10_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_11_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_11_Im; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_7; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_8; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_9; // @[FFTDesigns.scala 2750:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_10; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2750:28]
  wire [2:0] M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_8; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_9; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_10; // @[FFTDesigns.scala 2751:29]
  wire [3:0] M0_Config_ROM_io_out_11; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_8; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_9; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_10; // @[FFTDesigns.scala 2752:29]
  wire [3:0] M1_Config_ROM_io_out_11; // @[FFTDesigns.scala 2752:29]
  wire [2:0] Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2753:31]
  wire [3:0] Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2753:31]
  reg  offset_switch; // @[FFTDesigns.scala 2710:28]
  reg [2:0] cnt2; // @[FFTDesigns.scala 2755:25]
  reg [3:0] cnt; // @[FFTDesigns.scala 2756:24]
  wire [5:0] lo_lo = {io_in_en_5,io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2757:21]
  wire [11:0] lo = {io_in_en_11,io_in_en_10,io_in_en_9,io_in_en_8,io_in_en_7,io_in_en_6,lo_lo}; // @[FFTDesigns.scala 2757:21]
  wire [5:0] hi_lo = {io_in_en_17,io_in_en_16,io_in_en_15,io_in_en_14,io_in_en_13,io_in_en_12}; // @[FFTDesigns.scala 2757:21]
  wire [24:0] _T = {io_in_en_24,io_in_en_23,io_in_en_22,io_in_en_21,io_in_en_20,io_in_en_19,io_in_en_18,hi_lo,lo}; // @[FFTDesigns.scala 2757:21]
  wire  M0_0_re = |_T; // @[FFTDesigns.scala 2757:28]
  wire  _T_2 = cnt2 == 3'h7; // @[FFTDesigns.scala 2758:19]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2761:28]
  wire [3:0] _cnt_T_1 = cnt + 4'h1; // @[FFTDesigns.scala 2764:22]
  wire [2:0] _cnt2_T_1 = cnt2 + 3'h1; // @[FFTDesigns.scala 2767:24]
  wire  _GEN_5 = cnt2 == 3'h7 & cnt == 4'hb ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2758:69 2761:25]
  wire [4:0] _M0_0_in_raddr_T_1 = 4'h8 * _offset_switch_T; // @[FFTDesigns.scala 2778:56]
  wire [4:0] _GEN_862 = {{1'd0}, M0_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_0_in_raddr_T_3 = _GEN_862 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_863 = {{2'd0}, cnt2}; // @[FFTDesigns.scala 2781:34]
  wire [4:0] _M1_0_in_raddr_T_3 = _GEN_863 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2781:34]
  wire [4:0] _M1_0_in_waddr_T = 4'h8 * offset_switch; // @[FFTDesigns.scala 2782:56]
  wire [4:0] _GEN_864 = {{1'd0}, M1_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_0_in_waddr_T_2 = _GEN_864 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_865 = {{1'd0}, M0_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_1_in_raddr_T_3 = _GEN_865 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_867 = {{1'd0}, M1_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_1_in_waddr_T_2 = _GEN_867 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_868 = {{1'd0}, M0_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_2_in_raddr_T_3 = _GEN_868 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_870 = {{1'd0}, M1_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_2_in_waddr_T_2 = _GEN_870 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_871 = {{1'd0}, M0_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_3_in_raddr_T_3 = _GEN_871 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_873 = {{1'd0}, M1_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_3_in_waddr_T_2 = _GEN_873 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_874 = {{1'd0}, M0_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_4_in_raddr_T_3 = _GEN_874 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_876 = {{1'd0}, M1_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_4_in_waddr_T_2 = _GEN_876 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_877 = {{1'd0}, M0_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_5_in_raddr_T_3 = _GEN_877 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_879 = {{1'd0}, M1_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_5_in_waddr_T_2 = _GEN_879 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_880 = {{1'd0}, M0_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_6_in_raddr_T_3 = _GEN_880 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_882 = {{1'd0}, M1_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_6_in_waddr_T_2 = _GEN_882 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_883 = {{1'd0}, M0_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_7_in_raddr_T_3 = _GEN_883 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_885 = {{1'd0}, M1_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_7_in_waddr_T_2 = _GEN_885 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_886 = {{1'd0}, M0_Config_ROM_io_out_8}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_8_in_raddr_T_3 = _GEN_886 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_888 = {{1'd0}, M1_Config_ROM_io_out_8}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_8_in_waddr_T_2 = _GEN_888 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_889 = {{1'd0}, M0_Config_ROM_io_out_9}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_9_in_raddr_T_3 = _GEN_889 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_891 = {{1'd0}, M1_Config_ROM_io_out_9}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_9_in_waddr_T_2 = _GEN_891 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_892 = {{1'd0}, M0_Config_ROM_io_out_10}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_10_in_raddr_T_3 = _GEN_892 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_894 = {{1'd0}, M1_Config_ROM_io_out_10}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_10_in_waddr_T_2 = _GEN_894 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_895 = {{1'd0}, M0_Config_ROM_io_out_11}; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _M0_11_in_raddr_T_3 = _GEN_895 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [4:0] _GEN_897 = {{1'd0}, M1_Config_ROM_io_out_11}; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _M1_11_in_waddr_T_2 = _GEN_897 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [4:0] _GEN_7 = 4'h1 == cnt ? 5'h8 : 5'h0; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_8 = 4'h2 == cnt ? 5'h4 : _GEN_7; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_9 = 4'h3 == cnt ? 5'h0 : _GEN_8; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_10 = 4'h4 == cnt ? 5'h8 : _GEN_9; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_11 = 4'h5 == cnt ? 5'h4 : _GEN_10; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_12 = 4'h6 == cnt ? 5'h0 : _GEN_11; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_13 = 4'h7 == cnt ? 5'h8 : _GEN_12; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_14 = 4'h8 == cnt ? 5'h4 : _GEN_13; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_15 = 4'h9 == cnt ? 5'h0 : _GEN_14; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_16 = 4'ha == cnt ? 5'h8 : _GEN_15; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_17 = 4'hb == cnt ? 5'h4 : _GEN_16; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_20 = 4'h2 == cnt ? 5'h1 : 5'h0; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_21 = 4'h3 == cnt ? 5'h2 : _GEN_20; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_22 = 4'h4 == cnt ? 5'h2 : _GEN_21; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_23 = 4'h5 == cnt ? 5'h3 : _GEN_22; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_24 = 4'h6 == cnt ? 5'h4 : _GEN_23; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_25 = 4'h7 == cnt ? 5'h4 : _GEN_24; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_26 = 4'h8 == cnt ? 5'h5 : _GEN_25; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_27 = 4'h9 == cnt ? 5'h6 : _GEN_26; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_28 = 4'ha == cnt ? 5'h6 : _GEN_27; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_29 = 4'hb == cnt ? 5'h7 : _GEN_28; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _M0_0_in_waddr_T_2 = _GEN_29 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2799:50]
  wire [4:0] _GEN_31 = _GEN_17 == 5'h0 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_32 = _GEN_17 == 5'h0 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_33 = _GEN_17 == 5'h0 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_36 = 4'h1 == cnt ? 5'h9 : 5'h1; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_37 = 4'h2 == cnt ? 5'h5 : _GEN_36; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_38 = 4'h3 == cnt ? 5'h1 : _GEN_37; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_39 = 4'h4 == cnt ? 5'h9 : _GEN_38; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_40 = 4'h5 == cnt ? 5'h5 : _GEN_39; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_41 = 4'h6 == cnt ? 5'h1 : _GEN_40; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_42 = 4'h7 == cnt ? 5'h9 : _GEN_41; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_43 = 4'h8 == cnt ? 5'h5 : _GEN_42; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_44 = 4'h9 == cnt ? 5'h1 : _GEN_43; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_45 = 4'ha == cnt ? 5'h9 : _GEN_44; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_46 = 4'hb == cnt ? 5'h5 : _GEN_45; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_60 = _GEN_46 == 5'h0 ? _M0_0_in_waddr_T_2 : _GEN_31; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_61 = _GEN_46 == 5'h0 ? io_in_1_Im : _GEN_32; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_62 = _GEN_46 == 5'h0 ? io_in_1_Re : _GEN_33; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_65 = 4'h1 == cnt ? 5'ha : 5'h2; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_66 = 4'h2 == cnt ? 5'h6 : _GEN_65; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_67 = 4'h3 == cnt ? 5'h2 : _GEN_66; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_68 = 4'h4 == cnt ? 5'ha : _GEN_67; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_69 = 4'h5 == cnt ? 5'h6 : _GEN_68; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_70 = 4'h6 == cnt ? 5'h2 : _GEN_69; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_71 = 4'h7 == cnt ? 5'ha : _GEN_70; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_72 = 4'h8 == cnt ? 5'h6 : _GEN_71; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_73 = 4'h9 == cnt ? 5'h2 : _GEN_72; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_74 = 4'ha == cnt ? 5'ha : _GEN_73; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_75 = 4'hb == cnt ? 5'h6 : _GEN_74; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_89 = _GEN_75 == 5'h0 ? _M0_0_in_waddr_T_2 : _GEN_60; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_90 = _GEN_75 == 5'h0 ? io_in_2_Im : _GEN_61; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_91 = _GEN_75 == 5'h0 ? io_in_2_Re : _GEN_62; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_94 = 4'h1 == cnt ? 5'hb : 5'h3; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_95 = 4'h2 == cnt ? 5'h7 : _GEN_94; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_96 = 4'h3 == cnt ? 5'h3 : _GEN_95; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_97 = 4'h4 == cnt ? 5'hb : _GEN_96; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_98 = 4'h5 == cnt ? 5'h7 : _GEN_97; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_99 = 4'h6 == cnt ? 5'h3 : _GEN_98; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_100 = 4'h7 == cnt ? 5'hb : _GEN_99; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_101 = 4'h8 == cnt ? 5'h7 : _GEN_100; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_102 = 4'h9 == cnt ? 5'h3 : _GEN_101; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_103 = 4'ha == cnt ? 5'hb : _GEN_102; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_104 = 4'hb == cnt ? 5'h7 : _GEN_103; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_118 = _GEN_104 == 5'h0 ? _M0_0_in_waddr_T_2 : _GEN_89; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_119 = _GEN_104 == 5'h0 ? io_in_3_Im : _GEN_90; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_120 = _GEN_104 == 5'h0 ? io_in_3_Re : _GEN_91; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_123 = 4'h1 == cnt ? 5'h0 : 5'h4; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_124 = 4'h2 == cnt ? 5'h8 : _GEN_123; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_125 = 4'h3 == cnt ? 5'h4 : _GEN_124; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_126 = 4'h4 == cnt ? 5'h0 : _GEN_125; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_127 = 4'h5 == cnt ? 5'h8 : _GEN_126; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_128 = 4'h6 == cnt ? 5'h4 : _GEN_127; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_129 = 4'h7 == cnt ? 5'h0 : _GEN_128; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_130 = 4'h8 == cnt ? 5'h8 : _GEN_129; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_131 = 4'h9 == cnt ? 5'h4 : _GEN_130; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_132 = 4'ha == cnt ? 5'h0 : _GEN_131; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_133 = 4'hb == cnt ? 5'h8 : _GEN_132; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_135 = 4'h1 == cnt ? 5'h1 : 5'h0; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_136 = 4'h2 == cnt ? 5'h1 : _GEN_135; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_137 = 4'h3 == cnt ? 5'h2 : _GEN_136; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_138 = 4'h4 == cnt ? 5'h3 : _GEN_137; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_139 = 4'h5 == cnt ? 5'h3 : _GEN_138; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_140 = 4'h6 == cnt ? 5'h4 : _GEN_139; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_141 = 4'h7 == cnt ? 5'h5 : _GEN_140; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_142 = 4'h8 == cnt ? 5'h5 : _GEN_141; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_143 = 4'h9 == cnt ? 5'h6 : _GEN_142; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_144 = 4'ha == cnt ? 5'h7 : _GEN_143; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _GEN_145 = 4'hb == cnt ? 5'h7 : _GEN_144; // @[FFTDesigns.scala 2799:{50,50}]
  wire [4:0] _M0_0_in_waddr_T_14 = _GEN_145 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2799:50]
  wire [4:0] _GEN_147 = _GEN_133 == 5'h0 ? _M0_0_in_waddr_T_14 : _GEN_118; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_148 = _GEN_133 == 5'h0 ? io_in_4_Im : _GEN_119; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_149 = _GEN_133 == 5'h0 ? io_in_4_Re : _GEN_120; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_152 = 4'h1 == cnt ? 5'h1 : 5'h5; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_153 = 4'h2 == cnt ? 5'h9 : _GEN_152; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_154 = 4'h3 == cnt ? 5'h5 : _GEN_153; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_155 = 4'h4 == cnt ? 5'h1 : _GEN_154; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_156 = 4'h5 == cnt ? 5'h9 : _GEN_155; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_157 = 4'h6 == cnt ? 5'h5 : _GEN_156; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_158 = 4'h7 == cnt ? 5'h1 : _GEN_157; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_159 = 4'h8 == cnt ? 5'h9 : _GEN_158; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_160 = 4'h9 == cnt ? 5'h5 : _GEN_159; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_161 = 4'ha == cnt ? 5'h1 : _GEN_160; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_162 = 4'hb == cnt ? 5'h9 : _GEN_161; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_176 = _GEN_162 == 5'h0 ? _M0_0_in_waddr_T_14 : _GEN_147; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_177 = _GEN_162 == 5'h0 ? io_in_5_Im : _GEN_148; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_178 = _GEN_162 == 5'h0 ? io_in_5_Re : _GEN_149; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_181 = 4'h1 == cnt ? 5'h2 : 5'h6; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_182 = 4'h2 == cnt ? 5'ha : _GEN_181; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_183 = 4'h3 == cnt ? 5'h6 : _GEN_182; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_184 = 4'h4 == cnt ? 5'h2 : _GEN_183; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_185 = 4'h5 == cnt ? 5'ha : _GEN_184; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_186 = 4'h6 == cnt ? 5'h6 : _GEN_185; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_187 = 4'h7 == cnt ? 5'h2 : _GEN_186; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_188 = 4'h8 == cnt ? 5'ha : _GEN_187; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_189 = 4'h9 == cnt ? 5'h6 : _GEN_188; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_190 = 4'ha == cnt ? 5'h2 : _GEN_189; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_191 = 4'hb == cnt ? 5'ha : _GEN_190; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_205 = _GEN_191 == 5'h0 ? _M0_0_in_waddr_T_14 : _GEN_176; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_206 = _GEN_191 == 5'h0 ? io_in_6_Im : _GEN_177; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_207 = _GEN_191 == 5'h0 ? io_in_6_Re : _GEN_178; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_210 = 4'h1 == cnt ? 5'h3 : 5'h7; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_211 = 4'h2 == cnt ? 5'hb : _GEN_210; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_212 = 4'h3 == cnt ? 5'h7 : _GEN_211; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_213 = 4'h4 == cnt ? 5'h3 : _GEN_212; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_214 = 4'h5 == cnt ? 5'hb : _GEN_213; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_215 = 4'h6 == cnt ? 5'h7 : _GEN_214; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_216 = 4'h7 == cnt ? 5'h3 : _GEN_215; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_217 = 4'h8 == cnt ? 5'hb : _GEN_216; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_218 = 4'h9 == cnt ? 5'h7 : _GEN_217; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_219 = 4'ha == cnt ? 5'h3 : _GEN_218; // @[FFTDesigns.scala 2797:{35,35}]
  wire [4:0] _GEN_220 = 4'hb == cnt ? 5'hb : _GEN_219; // @[FFTDesigns.scala 2797:{35,35}]
  wire  _GEN_233 = _GEN_220 == 5'h0 | (_GEN_191 == 5'h0 | (_GEN_162 == 5'h0 | (_GEN_133 == 5'h0 | (_GEN_104 == 5'h0 | (
    _GEN_75 == 5'h0 | (_GEN_46 == 5'h0 | _GEN_17 == 5'h0)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_234 = _GEN_220 == 5'h0 ? _M0_0_in_waddr_T_14 : _GEN_205; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_235 = _GEN_220 == 5'h0 ? io_in_7_Im : _GEN_206; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_236 = _GEN_220 == 5'h0 ? io_in_7_Re : _GEN_207; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_239 = _GEN_17 == 5'h1 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_240 = _GEN_17 == 5'h1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_241 = _GEN_17 == 5'h1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_244 = _GEN_46 == 5'h1 ? _M0_0_in_waddr_T_2 : _GEN_239; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_245 = _GEN_46 == 5'h1 ? io_in_1_Im : _GEN_240; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_246 = _GEN_46 == 5'h1 ? io_in_1_Re : _GEN_241; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_249 = _GEN_75 == 5'h1 ? _M0_0_in_waddr_T_2 : _GEN_244; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_250 = _GEN_75 == 5'h1 ? io_in_2_Im : _GEN_245; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_251 = _GEN_75 == 5'h1 ? io_in_2_Re : _GEN_246; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_254 = _GEN_104 == 5'h1 ? _M0_0_in_waddr_T_2 : _GEN_249; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_255 = _GEN_104 == 5'h1 ? io_in_3_Im : _GEN_250; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_256 = _GEN_104 == 5'h1 ? io_in_3_Re : _GEN_251; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_259 = _GEN_133 == 5'h1 ? _M0_0_in_waddr_T_14 : _GEN_254; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_260 = _GEN_133 == 5'h1 ? io_in_4_Im : _GEN_255; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_261 = _GEN_133 == 5'h1 ? io_in_4_Re : _GEN_256; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_264 = _GEN_162 == 5'h1 ? _M0_0_in_waddr_T_14 : _GEN_259; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_265 = _GEN_162 == 5'h1 ? io_in_5_Im : _GEN_260; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_266 = _GEN_162 == 5'h1 ? io_in_5_Re : _GEN_261; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_269 = _GEN_191 == 5'h1 ? _M0_0_in_waddr_T_14 : _GEN_264; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_270 = _GEN_191 == 5'h1 ? io_in_6_Im : _GEN_265; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_271 = _GEN_191 == 5'h1 ? io_in_6_Re : _GEN_266; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_273 = _GEN_220 == 5'h1 | (_GEN_191 == 5'h1 | (_GEN_162 == 5'h1 | (_GEN_133 == 5'h1 | (_GEN_104 == 5'h1 | (
    _GEN_75 == 5'h1 | (_GEN_46 == 5'h1 | _GEN_17 == 5'h1)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_274 = _GEN_220 == 5'h1 ? _M0_0_in_waddr_T_14 : _GEN_269; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_275 = _GEN_220 == 5'h1 ? io_in_7_Im : _GEN_270; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_276 = _GEN_220 == 5'h1 ? io_in_7_Re : _GEN_271; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_279 = _GEN_17 == 5'h2 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_280 = _GEN_17 == 5'h2 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_281 = _GEN_17 == 5'h2 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_284 = _GEN_46 == 5'h2 ? _M0_0_in_waddr_T_2 : _GEN_279; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_285 = _GEN_46 == 5'h2 ? io_in_1_Im : _GEN_280; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_286 = _GEN_46 == 5'h2 ? io_in_1_Re : _GEN_281; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_289 = _GEN_75 == 5'h2 ? _M0_0_in_waddr_T_2 : _GEN_284; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_290 = _GEN_75 == 5'h2 ? io_in_2_Im : _GEN_285; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_291 = _GEN_75 == 5'h2 ? io_in_2_Re : _GEN_286; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_294 = _GEN_104 == 5'h2 ? _M0_0_in_waddr_T_2 : _GEN_289; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_295 = _GEN_104 == 5'h2 ? io_in_3_Im : _GEN_290; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_296 = _GEN_104 == 5'h2 ? io_in_3_Re : _GEN_291; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_299 = _GEN_133 == 5'h2 ? _M0_0_in_waddr_T_14 : _GEN_294; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_300 = _GEN_133 == 5'h2 ? io_in_4_Im : _GEN_295; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_301 = _GEN_133 == 5'h2 ? io_in_4_Re : _GEN_296; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_304 = _GEN_162 == 5'h2 ? _M0_0_in_waddr_T_14 : _GEN_299; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_305 = _GEN_162 == 5'h2 ? io_in_5_Im : _GEN_300; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_306 = _GEN_162 == 5'h2 ? io_in_5_Re : _GEN_301; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_309 = _GEN_191 == 5'h2 ? _M0_0_in_waddr_T_14 : _GEN_304; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_310 = _GEN_191 == 5'h2 ? io_in_6_Im : _GEN_305; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_311 = _GEN_191 == 5'h2 ? io_in_6_Re : _GEN_306; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_313 = _GEN_220 == 5'h2 | (_GEN_191 == 5'h2 | (_GEN_162 == 5'h2 | (_GEN_133 == 5'h2 | (_GEN_104 == 5'h2 | (
    _GEN_75 == 5'h2 | (_GEN_46 == 5'h2 | _GEN_17 == 5'h2)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_314 = _GEN_220 == 5'h2 ? _M0_0_in_waddr_T_14 : _GEN_309; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_315 = _GEN_220 == 5'h2 ? io_in_7_Im : _GEN_310; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_316 = _GEN_220 == 5'h2 ? io_in_7_Re : _GEN_311; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_319 = _GEN_17 == 5'h3 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_320 = _GEN_17 == 5'h3 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_321 = _GEN_17 == 5'h3 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_324 = _GEN_46 == 5'h3 ? _M0_0_in_waddr_T_2 : _GEN_319; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_325 = _GEN_46 == 5'h3 ? io_in_1_Im : _GEN_320; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_326 = _GEN_46 == 5'h3 ? io_in_1_Re : _GEN_321; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_329 = _GEN_75 == 5'h3 ? _M0_0_in_waddr_T_2 : _GEN_324; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_330 = _GEN_75 == 5'h3 ? io_in_2_Im : _GEN_325; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_331 = _GEN_75 == 5'h3 ? io_in_2_Re : _GEN_326; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_334 = _GEN_104 == 5'h3 ? _M0_0_in_waddr_T_2 : _GEN_329; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_335 = _GEN_104 == 5'h3 ? io_in_3_Im : _GEN_330; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_336 = _GEN_104 == 5'h3 ? io_in_3_Re : _GEN_331; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_339 = _GEN_133 == 5'h3 ? _M0_0_in_waddr_T_14 : _GEN_334; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_340 = _GEN_133 == 5'h3 ? io_in_4_Im : _GEN_335; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_341 = _GEN_133 == 5'h3 ? io_in_4_Re : _GEN_336; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_344 = _GEN_162 == 5'h3 ? _M0_0_in_waddr_T_14 : _GEN_339; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_345 = _GEN_162 == 5'h3 ? io_in_5_Im : _GEN_340; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_346 = _GEN_162 == 5'h3 ? io_in_5_Re : _GEN_341; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_349 = _GEN_191 == 5'h3 ? _M0_0_in_waddr_T_14 : _GEN_344; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_350 = _GEN_191 == 5'h3 ? io_in_6_Im : _GEN_345; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_351 = _GEN_191 == 5'h3 ? io_in_6_Re : _GEN_346; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_353 = _GEN_220 == 5'h3 | (_GEN_191 == 5'h3 | (_GEN_162 == 5'h3 | (_GEN_133 == 5'h3 | (_GEN_104 == 5'h3 | (
    _GEN_75 == 5'h3 | (_GEN_46 == 5'h3 | _GEN_17 == 5'h3)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_354 = _GEN_220 == 5'h3 ? _M0_0_in_waddr_T_14 : _GEN_349; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_355 = _GEN_220 == 5'h3 ? io_in_7_Im : _GEN_350; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_356 = _GEN_220 == 5'h3 ? io_in_7_Re : _GEN_351; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_359 = _GEN_17 == 5'h4 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_360 = _GEN_17 == 5'h4 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_361 = _GEN_17 == 5'h4 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_364 = _GEN_46 == 5'h4 ? _M0_0_in_waddr_T_2 : _GEN_359; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_365 = _GEN_46 == 5'h4 ? io_in_1_Im : _GEN_360; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_366 = _GEN_46 == 5'h4 ? io_in_1_Re : _GEN_361; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_369 = _GEN_75 == 5'h4 ? _M0_0_in_waddr_T_2 : _GEN_364; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_370 = _GEN_75 == 5'h4 ? io_in_2_Im : _GEN_365; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_371 = _GEN_75 == 5'h4 ? io_in_2_Re : _GEN_366; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_374 = _GEN_104 == 5'h4 ? _M0_0_in_waddr_T_2 : _GEN_369; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_375 = _GEN_104 == 5'h4 ? io_in_3_Im : _GEN_370; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_376 = _GEN_104 == 5'h4 ? io_in_3_Re : _GEN_371; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_379 = _GEN_133 == 5'h4 ? _M0_0_in_waddr_T_14 : _GEN_374; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_380 = _GEN_133 == 5'h4 ? io_in_4_Im : _GEN_375; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_381 = _GEN_133 == 5'h4 ? io_in_4_Re : _GEN_376; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_384 = _GEN_162 == 5'h4 ? _M0_0_in_waddr_T_14 : _GEN_379; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_385 = _GEN_162 == 5'h4 ? io_in_5_Im : _GEN_380; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_386 = _GEN_162 == 5'h4 ? io_in_5_Re : _GEN_381; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_389 = _GEN_191 == 5'h4 ? _M0_0_in_waddr_T_14 : _GEN_384; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_390 = _GEN_191 == 5'h4 ? io_in_6_Im : _GEN_385; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_391 = _GEN_191 == 5'h4 ? io_in_6_Re : _GEN_386; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_393 = _GEN_220 == 5'h4 | (_GEN_191 == 5'h4 | (_GEN_162 == 5'h4 | (_GEN_133 == 5'h4 | (_GEN_104 == 5'h4 | (
    _GEN_75 == 5'h4 | (_GEN_46 == 5'h4 | _GEN_17 == 5'h4)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_394 = _GEN_220 == 5'h4 ? _M0_0_in_waddr_T_14 : _GEN_389; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_395 = _GEN_220 == 5'h4 ? io_in_7_Im : _GEN_390; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_396 = _GEN_220 == 5'h4 ? io_in_7_Re : _GEN_391; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_399 = _GEN_17 == 5'h5 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_400 = _GEN_17 == 5'h5 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_401 = _GEN_17 == 5'h5 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_404 = _GEN_46 == 5'h5 ? _M0_0_in_waddr_T_2 : _GEN_399; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_405 = _GEN_46 == 5'h5 ? io_in_1_Im : _GEN_400; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_406 = _GEN_46 == 5'h5 ? io_in_1_Re : _GEN_401; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_409 = _GEN_75 == 5'h5 ? _M0_0_in_waddr_T_2 : _GEN_404; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_410 = _GEN_75 == 5'h5 ? io_in_2_Im : _GEN_405; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_411 = _GEN_75 == 5'h5 ? io_in_2_Re : _GEN_406; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_414 = _GEN_104 == 5'h5 ? _M0_0_in_waddr_T_2 : _GEN_409; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_415 = _GEN_104 == 5'h5 ? io_in_3_Im : _GEN_410; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_416 = _GEN_104 == 5'h5 ? io_in_3_Re : _GEN_411; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_419 = _GEN_133 == 5'h5 ? _M0_0_in_waddr_T_14 : _GEN_414; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_420 = _GEN_133 == 5'h5 ? io_in_4_Im : _GEN_415; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_421 = _GEN_133 == 5'h5 ? io_in_4_Re : _GEN_416; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_424 = _GEN_162 == 5'h5 ? _M0_0_in_waddr_T_14 : _GEN_419; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_425 = _GEN_162 == 5'h5 ? io_in_5_Im : _GEN_420; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_426 = _GEN_162 == 5'h5 ? io_in_5_Re : _GEN_421; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_429 = _GEN_191 == 5'h5 ? _M0_0_in_waddr_T_14 : _GEN_424; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_430 = _GEN_191 == 5'h5 ? io_in_6_Im : _GEN_425; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_431 = _GEN_191 == 5'h5 ? io_in_6_Re : _GEN_426; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_433 = _GEN_220 == 5'h5 | (_GEN_191 == 5'h5 | (_GEN_162 == 5'h5 | (_GEN_133 == 5'h5 | (_GEN_104 == 5'h5 | (
    _GEN_75 == 5'h5 | (_GEN_46 == 5'h5 | _GEN_17 == 5'h5)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_434 = _GEN_220 == 5'h5 ? _M0_0_in_waddr_T_14 : _GEN_429; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_435 = _GEN_220 == 5'h5 ? io_in_7_Im : _GEN_430; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_436 = _GEN_220 == 5'h5 ? io_in_7_Re : _GEN_431; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_439 = _GEN_17 == 5'h6 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_440 = _GEN_17 == 5'h6 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_441 = _GEN_17 == 5'h6 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_444 = _GEN_46 == 5'h6 ? _M0_0_in_waddr_T_2 : _GEN_439; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_445 = _GEN_46 == 5'h6 ? io_in_1_Im : _GEN_440; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_446 = _GEN_46 == 5'h6 ? io_in_1_Re : _GEN_441; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_449 = _GEN_75 == 5'h6 ? _M0_0_in_waddr_T_2 : _GEN_444; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_450 = _GEN_75 == 5'h6 ? io_in_2_Im : _GEN_445; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_451 = _GEN_75 == 5'h6 ? io_in_2_Re : _GEN_446; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_454 = _GEN_104 == 5'h6 ? _M0_0_in_waddr_T_2 : _GEN_449; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_455 = _GEN_104 == 5'h6 ? io_in_3_Im : _GEN_450; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_456 = _GEN_104 == 5'h6 ? io_in_3_Re : _GEN_451; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_459 = _GEN_133 == 5'h6 ? _M0_0_in_waddr_T_14 : _GEN_454; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_460 = _GEN_133 == 5'h6 ? io_in_4_Im : _GEN_455; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_461 = _GEN_133 == 5'h6 ? io_in_4_Re : _GEN_456; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_464 = _GEN_162 == 5'h6 ? _M0_0_in_waddr_T_14 : _GEN_459; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_465 = _GEN_162 == 5'h6 ? io_in_5_Im : _GEN_460; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_466 = _GEN_162 == 5'h6 ? io_in_5_Re : _GEN_461; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_469 = _GEN_191 == 5'h6 ? _M0_0_in_waddr_T_14 : _GEN_464; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_470 = _GEN_191 == 5'h6 ? io_in_6_Im : _GEN_465; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_471 = _GEN_191 == 5'h6 ? io_in_6_Re : _GEN_466; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_473 = _GEN_220 == 5'h6 | (_GEN_191 == 5'h6 | (_GEN_162 == 5'h6 | (_GEN_133 == 5'h6 | (_GEN_104 == 5'h6 | (
    _GEN_75 == 5'h6 | (_GEN_46 == 5'h6 | _GEN_17 == 5'h6)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_474 = _GEN_220 == 5'h6 ? _M0_0_in_waddr_T_14 : _GEN_469; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_475 = _GEN_220 == 5'h6 ? io_in_7_Im : _GEN_470; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_476 = _GEN_220 == 5'h6 ? io_in_7_Re : _GEN_471; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_479 = _GEN_17 == 5'h7 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_480 = _GEN_17 == 5'h7 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_481 = _GEN_17 == 5'h7 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_484 = _GEN_46 == 5'h7 ? _M0_0_in_waddr_T_2 : _GEN_479; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_485 = _GEN_46 == 5'h7 ? io_in_1_Im : _GEN_480; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_486 = _GEN_46 == 5'h7 ? io_in_1_Re : _GEN_481; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_489 = _GEN_75 == 5'h7 ? _M0_0_in_waddr_T_2 : _GEN_484; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_490 = _GEN_75 == 5'h7 ? io_in_2_Im : _GEN_485; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_491 = _GEN_75 == 5'h7 ? io_in_2_Re : _GEN_486; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_494 = _GEN_104 == 5'h7 ? _M0_0_in_waddr_T_2 : _GEN_489; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_495 = _GEN_104 == 5'h7 ? io_in_3_Im : _GEN_490; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_496 = _GEN_104 == 5'h7 ? io_in_3_Re : _GEN_491; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_499 = _GEN_133 == 5'h7 ? _M0_0_in_waddr_T_14 : _GEN_494; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_500 = _GEN_133 == 5'h7 ? io_in_4_Im : _GEN_495; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_501 = _GEN_133 == 5'h7 ? io_in_4_Re : _GEN_496; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_504 = _GEN_162 == 5'h7 ? _M0_0_in_waddr_T_14 : _GEN_499; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_505 = _GEN_162 == 5'h7 ? io_in_5_Im : _GEN_500; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_506 = _GEN_162 == 5'h7 ? io_in_5_Re : _GEN_501; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_509 = _GEN_191 == 5'h7 ? _M0_0_in_waddr_T_14 : _GEN_504; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_510 = _GEN_191 == 5'h7 ? io_in_6_Im : _GEN_505; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_511 = _GEN_191 == 5'h7 ? io_in_6_Re : _GEN_506; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_513 = _GEN_220 == 5'h7 | (_GEN_191 == 5'h7 | (_GEN_162 == 5'h7 | (_GEN_133 == 5'h7 | (_GEN_104 == 5'h7 | (
    _GEN_75 == 5'h7 | (_GEN_46 == 5'h7 | _GEN_17 == 5'h7)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_514 = _GEN_220 == 5'h7 ? _M0_0_in_waddr_T_14 : _GEN_509; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_515 = _GEN_220 == 5'h7 ? io_in_7_Im : _GEN_510; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_516 = _GEN_220 == 5'h7 ? io_in_7_Re : _GEN_511; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_519 = _GEN_17 == 5'h8 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_520 = _GEN_17 == 5'h8 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_521 = _GEN_17 == 5'h8 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_524 = _GEN_46 == 5'h8 ? _M0_0_in_waddr_T_2 : _GEN_519; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_525 = _GEN_46 == 5'h8 ? io_in_1_Im : _GEN_520; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_526 = _GEN_46 == 5'h8 ? io_in_1_Re : _GEN_521; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_529 = _GEN_75 == 5'h8 ? _M0_0_in_waddr_T_2 : _GEN_524; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_530 = _GEN_75 == 5'h8 ? io_in_2_Im : _GEN_525; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_531 = _GEN_75 == 5'h8 ? io_in_2_Re : _GEN_526; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_534 = _GEN_104 == 5'h8 ? _M0_0_in_waddr_T_2 : _GEN_529; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_535 = _GEN_104 == 5'h8 ? io_in_3_Im : _GEN_530; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_536 = _GEN_104 == 5'h8 ? io_in_3_Re : _GEN_531; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_539 = _GEN_133 == 5'h8 ? _M0_0_in_waddr_T_14 : _GEN_534; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_540 = _GEN_133 == 5'h8 ? io_in_4_Im : _GEN_535; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_541 = _GEN_133 == 5'h8 ? io_in_4_Re : _GEN_536; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_544 = _GEN_162 == 5'h8 ? _M0_0_in_waddr_T_14 : _GEN_539; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_545 = _GEN_162 == 5'h8 ? io_in_5_Im : _GEN_540; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_546 = _GEN_162 == 5'h8 ? io_in_5_Re : _GEN_541; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_549 = _GEN_191 == 5'h8 ? _M0_0_in_waddr_T_14 : _GEN_544; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_550 = _GEN_191 == 5'h8 ? io_in_6_Im : _GEN_545; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_551 = _GEN_191 == 5'h8 ? io_in_6_Re : _GEN_546; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_553 = _GEN_220 == 5'h8 | (_GEN_191 == 5'h8 | (_GEN_162 == 5'h8 | (_GEN_133 == 5'h8 | (_GEN_104 == 5'h8 | (
    _GEN_75 == 5'h8 | (_GEN_46 == 5'h8 | _GEN_17 == 5'h8)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_554 = _GEN_220 == 5'h8 ? _M0_0_in_waddr_T_14 : _GEN_549; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_555 = _GEN_220 == 5'h8 ? io_in_7_Im : _GEN_550; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_556 = _GEN_220 == 5'h8 ? io_in_7_Re : _GEN_551; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_559 = _GEN_17 == 5'h9 ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_560 = _GEN_17 == 5'h9 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_561 = _GEN_17 == 5'h9 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_564 = _GEN_46 == 5'h9 ? _M0_0_in_waddr_T_2 : _GEN_559; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_565 = _GEN_46 == 5'h9 ? io_in_1_Im : _GEN_560; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_566 = _GEN_46 == 5'h9 ? io_in_1_Re : _GEN_561; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_569 = _GEN_75 == 5'h9 ? _M0_0_in_waddr_T_2 : _GEN_564; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_570 = _GEN_75 == 5'h9 ? io_in_2_Im : _GEN_565; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_571 = _GEN_75 == 5'h9 ? io_in_2_Re : _GEN_566; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_574 = _GEN_104 == 5'h9 ? _M0_0_in_waddr_T_2 : _GEN_569; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_575 = _GEN_104 == 5'h9 ? io_in_3_Im : _GEN_570; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_576 = _GEN_104 == 5'h9 ? io_in_3_Re : _GEN_571; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_579 = _GEN_133 == 5'h9 ? _M0_0_in_waddr_T_14 : _GEN_574; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_580 = _GEN_133 == 5'h9 ? io_in_4_Im : _GEN_575; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_581 = _GEN_133 == 5'h9 ? io_in_4_Re : _GEN_576; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_584 = _GEN_162 == 5'h9 ? _M0_0_in_waddr_T_14 : _GEN_579; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_585 = _GEN_162 == 5'h9 ? io_in_5_Im : _GEN_580; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_586 = _GEN_162 == 5'h9 ? io_in_5_Re : _GEN_581; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_589 = _GEN_191 == 5'h9 ? _M0_0_in_waddr_T_14 : _GEN_584; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_590 = _GEN_191 == 5'h9 ? io_in_6_Im : _GEN_585; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_591 = _GEN_191 == 5'h9 ? io_in_6_Re : _GEN_586; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_593 = _GEN_220 == 5'h9 | (_GEN_191 == 5'h9 | (_GEN_162 == 5'h9 | (_GEN_133 == 5'h9 | (_GEN_104 == 5'h9 | (
    _GEN_75 == 5'h9 | (_GEN_46 == 5'h9 | _GEN_17 == 5'h9)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_594 = _GEN_220 == 5'h9 ? _M0_0_in_waddr_T_14 : _GEN_589; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_595 = _GEN_220 == 5'h9 ? io_in_7_Im : _GEN_590; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_596 = _GEN_220 == 5'h9 ? io_in_7_Re : _GEN_591; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_599 = _GEN_17 == 5'ha ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_600 = _GEN_17 == 5'ha ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_601 = _GEN_17 == 5'ha ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_604 = _GEN_46 == 5'ha ? _M0_0_in_waddr_T_2 : _GEN_599; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_605 = _GEN_46 == 5'ha ? io_in_1_Im : _GEN_600; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_606 = _GEN_46 == 5'ha ? io_in_1_Re : _GEN_601; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_609 = _GEN_75 == 5'ha ? _M0_0_in_waddr_T_2 : _GEN_604; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_610 = _GEN_75 == 5'ha ? io_in_2_Im : _GEN_605; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_611 = _GEN_75 == 5'ha ? io_in_2_Re : _GEN_606; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_614 = _GEN_104 == 5'ha ? _M0_0_in_waddr_T_2 : _GEN_609; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_615 = _GEN_104 == 5'ha ? io_in_3_Im : _GEN_610; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_616 = _GEN_104 == 5'ha ? io_in_3_Re : _GEN_611; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_619 = _GEN_133 == 5'ha ? _M0_0_in_waddr_T_14 : _GEN_614; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_620 = _GEN_133 == 5'ha ? io_in_4_Im : _GEN_615; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_621 = _GEN_133 == 5'ha ? io_in_4_Re : _GEN_616; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_624 = _GEN_162 == 5'ha ? _M0_0_in_waddr_T_14 : _GEN_619; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_625 = _GEN_162 == 5'ha ? io_in_5_Im : _GEN_620; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_626 = _GEN_162 == 5'ha ? io_in_5_Re : _GEN_621; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_629 = _GEN_191 == 5'ha ? _M0_0_in_waddr_T_14 : _GEN_624; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_630 = _GEN_191 == 5'ha ? io_in_6_Im : _GEN_625; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_631 = _GEN_191 == 5'ha ? io_in_6_Re : _GEN_626; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_633 = _GEN_220 == 5'ha | (_GEN_191 == 5'ha | (_GEN_162 == 5'ha | (_GEN_133 == 5'ha | (_GEN_104 == 5'ha | (
    _GEN_75 == 5'ha | (_GEN_46 == 5'ha | _GEN_17 == 5'ha)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_634 = _GEN_220 == 5'ha ? _M0_0_in_waddr_T_14 : _GEN_629; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_635 = _GEN_220 == 5'ha ? io_in_7_Im : _GEN_630; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_636 = _GEN_220 == 5'ha ? io_in_7_Re : _GEN_631; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_639 = _GEN_17 == 5'hb ? _M0_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_640 = _GEN_17 == 5'hb ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_641 = _GEN_17 == 5'hb ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [4:0] _GEN_644 = _GEN_46 == 5'hb ? _M0_0_in_waddr_T_2 : _GEN_639; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_645 = _GEN_46 == 5'hb ? io_in_1_Im : _GEN_640; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_646 = _GEN_46 == 5'hb ? io_in_1_Re : _GEN_641; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_649 = _GEN_75 == 5'hb ? _M0_0_in_waddr_T_2 : _GEN_644; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_650 = _GEN_75 == 5'hb ? io_in_2_Im : _GEN_645; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_651 = _GEN_75 == 5'hb ? io_in_2_Re : _GEN_646; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_654 = _GEN_104 == 5'hb ? _M0_0_in_waddr_T_2 : _GEN_649; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_655 = _GEN_104 == 5'hb ? io_in_3_Im : _GEN_650; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_656 = _GEN_104 == 5'hb ? io_in_3_Re : _GEN_651; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_659 = _GEN_133 == 5'hb ? _M0_0_in_waddr_T_14 : _GEN_654; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_660 = _GEN_133 == 5'hb ? io_in_4_Im : _GEN_655; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_661 = _GEN_133 == 5'hb ? io_in_4_Re : _GEN_656; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_664 = _GEN_162 == 5'hb ? _M0_0_in_waddr_T_14 : _GEN_659; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_665 = _GEN_162 == 5'hb ? io_in_5_Im : _GEN_660; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_666 = _GEN_162 == 5'hb ? io_in_5_Re : _GEN_661; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_669 = _GEN_191 == 5'hb ? _M0_0_in_waddr_T_14 : _GEN_664; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_670 = _GEN_191 == 5'hb ? io_in_6_Im : _GEN_665; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_671 = _GEN_191 == 5'hb ? io_in_6_Re : _GEN_666; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_673 = _GEN_220 == 5'hb | (_GEN_191 == 5'hb | (_GEN_162 == 5'hb | (_GEN_133 == 5'hb | (_GEN_104 == 5'hb | (
    _GEN_75 == 5'hb | (_GEN_46 == 5'hb | _GEN_17 == 5'hb)))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [4:0] _GEN_674 = _GEN_220 == 5'hb ? _M0_0_in_waddr_T_14 : _GEN_669; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_675 = _GEN_220 == 5'hb ? io_in_7_Im : _GEN_670; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_676 = _GEN_220 == 5'hb ? io_in_7_Re : _GEN_671; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [4:0] _GEN_682 = M0_0_re ? _M0_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_683 = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2781:26 2816:26]
  wire [4:0] _GEN_684 = M0_0_re ? _M1_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_692 = M0_0_re ? _M0_1_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_694 = M0_0_re ? _M1_1_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_702 = M0_0_re ? _M0_2_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_704 = M0_0_re ? _M1_2_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_712 = M0_0_re ? _M0_3_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_714 = M0_0_re ? _M1_3_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_722 = M0_0_re ? _M0_4_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_724 = M0_0_re ? _M1_4_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_732 = M0_0_re ? _M0_5_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_734 = M0_0_re ? _M1_5_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_742 = M0_0_re ? _M0_6_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_744 = M0_0_re ? _M1_6_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_752 = M0_0_re ? _M0_7_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_754 = M0_0_re ? _M1_7_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_762 = M0_0_re ? _M0_8_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_764 = M0_0_re ? _M1_8_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_772 = M0_0_re ? _M0_9_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_774 = M0_0_re ? _M1_9_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_782 = M0_0_re ? _M0_10_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_784 = M0_0_re ? _M1_10_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_792 = M0_0_re ? _M0_11_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [4:0] _GEN_794 = M0_0_re ? _M1_11_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [4:0] _GEN_803 = M0_0_re ? _GEN_234 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_808 = M0_0_re ? _GEN_274 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_813 = M0_0_re ? _GEN_314 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_818 = M0_0_re ? _GEN_354 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_823 = M0_0_re ? _GEN_394 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_828 = M0_0_re ? _GEN_434 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_833 = M0_0_re ? _GEN_474 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_838 = M0_0_re ? _GEN_514 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_843 = M0_0_re ? _GEN_554 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_848 = M0_0_re ? _GEN_594 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_853 = M0_0_re ? _GEN_634 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [4:0] _GEN_858 = M0_0_re ? _GEN_674 : 5'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  RAM_Block_112 RAM_Block ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_1 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_2 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_3 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_4 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_5 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_6 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_7 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_8 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_9 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_10 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_11 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_12 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_13 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_14 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_15 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_16 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_16_clock),
    .io_in_raddr(RAM_Block_16_io_in_raddr),
    .io_in_waddr(RAM_Block_16_io_in_waddr),
    .io_in_data_Re(RAM_Block_16_io_in_data_Re),
    .io_in_data_Im(RAM_Block_16_io_in_data_Im),
    .io_re(RAM_Block_16_io_re),
    .io_wr(RAM_Block_16_io_wr),
    .io_en(RAM_Block_16_io_en),
    .io_out_data_Re(RAM_Block_16_io_out_data_Re),
    .io_out_data_Im(RAM_Block_16_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_17 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_17_clock),
    .io_in_raddr(RAM_Block_17_io_in_raddr),
    .io_in_waddr(RAM_Block_17_io_in_waddr),
    .io_in_data_Re(RAM_Block_17_io_in_data_Re),
    .io_in_data_Im(RAM_Block_17_io_in_data_Im),
    .io_re(RAM_Block_17_io_re),
    .io_wr(RAM_Block_17_io_wr),
    .io_en(RAM_Block_17_io_en),
    .io_out_data_Re(RAM_Block_17_io_out_data_Re),
    .io_out_data_Im(RAM_Block_17_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_18 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_18_clock),
    .io_in_raddr(RAM_Block_18_io_in_raddr),
    .io_in_waddr(RAM_Block_18_io_in_waddr),
    .io_in_data_Re(RAM_Block_18_io_in_data_Re),
    .io_in_data_Im(RAM_Block_18_io_in_data_Im),
    .io_re(RAM_Block_18_io_re),
    .io_wr(RAM_Block_18_io_wr),
    .io_en(RAM_Block_18_io_en),
    .io_out_data_Re(RAM_Block_18_io_out_data_Re),
    .io_out_data_Im(RAM_Block_18_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_19 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_19_clock),
    .io_in_raddr(RAM_Block_19_io_in_raddr),
    .io_in_waddr(RAM_Block_19_io_in_waddr),
    .io_in_data_Re(RAM_Block_19_io_in_data_Re),
    .io_in_data_Im(RAM_Block_19_io_in_data_Im),
    .io_re(RAM_Block_19_io_re),
    .io_wr(RAM_Block_19_io_wr),
    .io_en(RAM_Block_19_io_en),
    .io_out_data_Re(RAM_Block_19_io_out_data_Re),
    .io_out_data_Im(RAM_Block_19_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_20 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_20_clock),
    .io_in_raddr(RAM_Block_20_io_in_raddr),
    .io_in_waddr(RAM_Block_20_io_in_waddr),
    .io_in_data_Re(RAM_Block_20_io_in_data_Re),
    .io_in_data_Im(RAM_Block_20_io_in_data_Im),
    .io_re(RAM_Block_20_io_re),
    .io_wr(RAM_Block_20_io_wr),
    .io_en(RAM_Block_20_io_en),
    .io_out_data_Re(RAM_Block_20_io_out_data_Re),
    .io_out_data_Im(RAM_Block_20_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_21 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_21_clock),
    .io_in_raddr(RAM_Block_21_io_in_raddr),
    .io_in_waddr(RAM_Block_21_io_in_waddr),
    .io_in_data_Re(RAM_Block_21_io_in_data_Re),
    .io_in_data_Im(RAM_Block_21_io_in_data_Im),
    .io_re(RAM_Block_21_io_re),
    .io_wr(RAM_Block_21_io_wr),
    .io_en(RAM_Block_21_io_en),
    .io_out_data_Re(RAM_Block_21_io_out_data_Re),
    .io_out_data_Im(RAM_Block_21_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_22 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_22_clock),
    .io_in_raddr(RAM_Block_22_io_in_raddr),
    .io_in_waddr(RAM_Block_22_io_in_waddr),
    .io_in_data_Re(RAM_Block_22_io_in_data_Re),
    .io_in_data_Im(RAM_Block_22_io_in_data_Im),
    .io_re(RAM_Block_22_io_re),
    .io_wr(RAM_Block_22_io_wr),
    .io_en(RAM_Block_22_io_en),
    .io_out_data_Re(RAM_Block_22_io_out_data_Re),
    .io_out_data_Im(RAM_Block_22_io_out_data_Im)
  );
  RAM_Block_112 RAM_Block_23 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_23_clock),
    .io_in_raddr(RAM_Block_23_io_in_raddr),
    .io_in_waddr(RAM_Block_23_io_in_waddr),
    .io_in_data_Re(RAM_Block_23_io_in_data_Re),
    .io_in_data_Im(RAM_Block_23_io_in_data_Im),
    .io_re(RAM_Block_23_io_re),
    .io_wr(RAM_Block_23_io_wr),
    .io_en(RAM_Block_23_io_en),
    .io_out_data_Re(RAM_Block_23_io_out_data_Re),
    .io_out_data_Im(RAM_Block_23_io_out_data_Im)
  );
  PermutationModuleStreamed_7 PermutationModuleStreamed ( // @[FFTDesigns.scala 2750:28]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_8_Re(PermutationModuleStreamed_io_in_8_Re),
    .io_in_8_Im(PermutationModuleStreamed_io_in_8_Im),
    .io_in_9_Re(PermutationModuleStreamed_io_in_9_Re),
    .io_in_9_Im(PermutationModuleStreamed_io_in_9_Im),
    .io_in_10_Re(PermutationModuleStreamed_io_in_10_Re),
    .io_in_10_Im(PermutationModuleStreamed_io_in_10_Im),
    .io_in_11_Re(PermutationModuleStreamed_io_in_11_Re),
    .io_in_11_Im(PermutationModuleStreamed_io_in_11_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_in_config_7(PermutationModuleStreamed_io_in_config_7),
    .io_in_config_8(PermutationModuleStreamed_io_in_config_8),
    .io_in_config_9(PermutationModuleStreamed_io_in_config_9),
    .io_in_config_10(PermutationModuleStreamed_io_in_config_10),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im),
    .io_out_8_Re(PermutationModuleStreamed_io_out_8_Re),
    .io_out_8_Im(PermutationModuleStreamed_io_out_8_Im),
    .io_out_9_Re(PermutationModuleStreamed_io_out_9_Re),
    .io_out_9_Im(PermutationModuleStreamed_io_out_9_Im),
    .io_out_10_Re(PermutationModuleStreamed_io_out_10_Re),
    .io_out_10_Im(PermutationModuleStreamed_io_out_10_Im),
    .io_out_11_Re(PermutationModuleStreamed_io_out_11_Re),
    .io_out_11_Im(PermutationModuleStreamed_io_out_11_Im)
  );
  M0_Config_ROM_7 M0_Config_ROM ( // @[FFTDesigns.scala 2751:29]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7),
    .io_out_8(M0_Config_ROM_io_out_8),
    .io_out_9(M0_Config_ROM_io_out_9),
    .io_out_10(M0_Config_ROM_io_out_10),
    .io_out_11(M0_Config_ROM_io_out_11)
  );
  M1_Config_ROM_7 M1_Config_ROM ( // @[FFTDesigns.scala 2752:29]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7),
    .io_out_8(M1_Config_ROM_io_out_8),
    .io_out_9(M1_Config_ROM_io_out_9),
    .io_out_10(M1_Config_ROM_io_out_10),
    .io_out_11(M1_Config_ROM_io_out_11)
  );
  Streaming_Permute_Config_7 Streaming_Permute_Config ( // @[FFTDesigns.scala 2753:31]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6),
    .io_out_7(Streaming_Permute_Config_io_out_7),
    .io_out_8(Streaming_Permute_Config_io_out_8),
    .io_out_9(Streaming_Permute_Config_io_out_9),
    .io_out_10(Streaming_Permute_Config_io_out_10)
  );
  assign io_out_0_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_0_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_1_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_1_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_2_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_2_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_3_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_3_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_4_Re = RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_4_Im = RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_5_Re = RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_5_Im = RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_6_Re = RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_6_Im = RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_7_Re = RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_7_Im = RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_8_Re = RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_8_Im = RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_9_Re = RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_9_Im = RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_10_Re = RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_10_Im = RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_11_Re = RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_11_Im = RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = _GEN_682[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_io_in_waddr = _GEN_803[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_io_in_data_Re = M0_0_re ? _GEN_236 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_io_in_data_Im = M0_0_re ? _GEN_235 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_io_wr = M0_0_re & _GEN_233; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = _GEN_692[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_1_io_in_waddr = _GEN_808[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_1_io_in_data_Re = M0_0_re ? _GEN_276 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_1_io_in_data_Im = M0_0_re ? _GEN_275 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_1_io_wr = M0_0_re & _GEN_273; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = _GEN_702[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_2_io_in_waddr = _GEN_813[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_2_io_in_data_Re = M0_0_re ? _GEN_316 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_2_io_in_data_Im = M0_0_re ? _GEN_315 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_2_io_wr = M0_0_re & _GEN_313; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = _GEN_712[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_3_io_in_waddr = _GEN_818[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_3_io_in_data_Re = M0_0_re ? _GEN_356 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_3_io_in_data_Im = M0_0_re ? _GEN_355 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_3_io_wr = M0_0_re & _GEN_353; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = _GEN_722[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_4_io_in_waddr = _GEN_823[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_4_io_in_data_Re = M0_0_re ? _GEN_396 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_4_io_in_data_Im = M0_0_re ? _GEN_395 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_4_io_wr = M0_0_re & _GEN_393; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = _GEN_732[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_5_io_in_waddr = _GEN_828[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_5_io_in_data_Re = M0_0_re ? _GEN_436 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_5_io_in_data_Im = M0_0_re ? _GEN_435 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_5_io_wr = M0_0_re & _GEN_433; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = _GEN_742[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_6_io_in_waddr = _GEN_833[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_6_io_in_data_Re = M0_0_re ? _GEN_476 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_6_io_in_data_Im = M0_0_re ? _GEN_475 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_6_io_wr = M0_0_re & _GEN_473; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = _GEN_752[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_7_io_in_waddr = _GEN_838[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_7_io_in_data_Re = M0_0_re ? _GEN_516 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_7_io_in_data_Im = M0_0_re ? _GEN_515 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_7_io_wr = M0_0_re & _GEN_513; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = _GEN_762[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_8_io_in_waddr = _GEN_843[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_8_io_in_data_Re = M0_0_re ? _GEN_556 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_8_io_in_data_Im = M0_0_re ? _GEN_555 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_8_io_wr = M0_0_re & _GEN_553; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = _GEN_772[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_9_io_in_waddr = _GEN_848[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_9_io_in_data_Re = M0_0_re ? _GEN_596 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_9_io_in_data_Im = M0_0_re ? _GEN_595 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_9_io_wr = M0_0_re & _GEN_593; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = _GEN_782[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_10_io_in_waddr = _GEN_853[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_10_io_in_data_Re = M0_0_re ? _GEN_636 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_10_io_in_data_Im = M0_0_re ? _GEN_635 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_10_io_wr = M0_0_re & _GEN_633; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = _GEN_792[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_11_io_in_waddr = _GEN_858[3:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_11_io_in_data_Re = M0_0_re ? _GEN_676 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_11_io_in_data_Im = M0_0_re ? _GEN_675 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_11_io_wr = M0_0_re & _GEN_673; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_12_io_in_waddr = _GEN_684[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_12_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_12_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_12_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_13_io_in_waddr = _GEN_694[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_13_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_13_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_13_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_14_io_in_waddr = _GEN_704[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_14_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_14_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_14_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_15_io_in_waddr = _GEN_714[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_15_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_15_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_15_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_16_clock = clock;
  assign RAM_Block_16_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_16_io_in_waddr = _GEN_724[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_16_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_16_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_16_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_16_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_16_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_17_clock = clock;
  assign RAM_Block_17_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_17_io_in_waddr = _GEN_734[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_17_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_17_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_17_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_17_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_17_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_18_clock = clock;
  assign RAM_Block_18_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_18_io_in_waddr = _GEN_744[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_18_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_18_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_18_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_18_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_18_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_19_clock = clock;
  assign RAM_Block_19_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_19_io_in_waddr = _GEN_754[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_19_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_19_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_19_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_19_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_19_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_20_clock = clock;
  assign RAM_Block_20_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_20_io_in_waddr = _GEN_764[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_20_io_in_data_Re = PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_20_io_in_data_Im = PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_20_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_20_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_20_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_21_clock = clock;
  assign RAM_Block_21_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_21_io_in_waddr = _GEN_774[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_21_io_in_data_Re = PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_21_io_in_data_Im = PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_21_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_21_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_21_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_22_clock = clock;
  assign RAM_Block_22_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_22_io_in_waddr = _GEN_784[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_22_io_in_data_Re = PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_22_io_in_data_Im = PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_22_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_22_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_22_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_23_clock = clock;
  assign RAM_Block_23_io_in_raddr = _GEN_683[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_23_io_in_waddr = _GEN_794[3:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_23_io_in_data_Re = PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_23_io_in_data_Im = PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_23_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_23_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_23_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_8_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_8_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_9_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_9_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_10_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_10_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_11_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_11_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_7 = Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_8 = Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_9 = Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_10 = Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign M0_Config_ROM_io_in_cnt = cnt2; // @[FFTDesigns.scala 2829:24]
  assign M1_Config_ROM_io_in_cnt = cnt2; // @[FFTDesigns.scala 2830:24]
  assign Streaming_Permute_Config_io_in_cnt = cnt2; // @[FFTDesigns.scala 2831:26]
  always @(posedge clock) begin
    offset_switch <= M0_0_re & _GEN_5; // @[FFTDesigns.scala 2757:33 2825:23]
    if (reset) begin // @[FFTDesigns.scala 2755:25]
      cnt2 <= 3'h0; // @[FFTDesigns.scala 2755:25]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2757:33]
      if (cnt2 == 3'h7 & cnt == 4'hb) begin // @[FFTDesigns.scala 2758:69]
        cnt2 <= 3'h0; // @[FFTDesigns.scala 2759:16]
      end else if (!(_T_2)) begin // @[FFTDesigns.scala 2762:46]
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2767:16]
      end
    end
    if (reset) begin // @[FFTDesigns.scala 2756:24]
      cnt <= 4'h0; // @[FFTDesigns.scala 2756:24]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2757:33]
      if (cnt2 == 3'h7 & cnt == 4'hb) begin // @[FFTDesigns.scala 2758:69]
        cnt <= 4'h0; // @[FFTDesigns.scala 2760:15]
      end else if (_T_2) begin // @[FFTDesigns.scala 2762:46]
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2764:15]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2768:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt2 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  cnt = _RAND_2[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_Block_mw(
  input         clock,
  input  [4:0]  io_in_raddr,
  input  [4:0]  io_in_waddr_0,
  input  [4:0]  io_in_waddr_1,
  input  [31:0] io_in_data_0_Re,
  input  [31:0] io_in_data_0_Im,
  input  [31:0] io_in_data_1_Re,
  input  [31:0] io_in_data_1_Im,
  input         io_re,
  input         io_wr_0,
  input         io_wr_1,
  input         io_en,
  output [31:0] io_out_data_Re,
  output [31:0] io_out_data_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_0_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_1_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_1_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_2_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_2_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_3_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_3_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_4_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_4_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_5_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_5_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_6_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_6_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_7_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_7_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_8_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_8_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_9_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_9_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_10_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_10_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_11_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_11_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_12_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_12_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_13_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_13_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_14_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_14_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_15_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_15_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_16_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_16_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_17_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_17_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_18_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_18_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_19_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_19_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_20_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_20_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_21_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_21_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_22_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_22_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_23_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_23_Im; // @[FFTDesigns.scala 3313:18]
  wire [31:0] _GEN_0 = 5'h0 == io_in_waddr_0 ? io_in_data_0_Im : mem_0_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_1 = 5'h1 == io_in_waddr_0 ? io_in_data_0_Im : mem_1_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_2 = 5'h2 == io_in_waddr_0 ? io_in_data_0_Im : mem_2_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_3 = 5'h3 == io_in_waddr_0 ? io_in_data_0_Im : mem_3_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_4 = 5'h4 == io_in_waddr_0 ? io_in_data_0_Im : mem_4_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_5 = 5'h5 == io_in_waddr_0 ? io_in_data_0_Im : mem_5_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_6 = 5'h6 == io_in_waddr_0 ? io_in_data_0_Im : mem_6_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_7 = 5'h7 == io_in_waddr_0 ? io_in_data_0_Im : mem_7_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_8 = 5'h8 == io_in_waddr_0 ? io_in_data_0_Im : mem_8_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_9 = 5'h9 == io_in_waddr_0 ? io_in_data_0_Im : mem_9_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_10 = 5'ha == io_in_waddr_0 ? io_in_data_0_Im : mem_10_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_11 = 5'hb == io_in_waddr_0 ? io_in_data_0_Im : mem_11_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_12 = 5'hc == io_in_waddr_0 ? io_in_data_0_Im : mem_12_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_13 = 5'hd == io_in_waddr_0 ? io_in_data_0_Im : mem_13_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_14 = 5'he == io_in_waddr_0 ? io_in_data_0_Im : mem_14_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_15 = 5'hf == io_in_waddr_0 ? io_in_data_0_Im : mem_15_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_16 = 5'h10 == io_in_waddr_0 ? io_in_data_0_Im : mem_16_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_17 = 5'h11 == io_in_waddr_0 ? io_in_data_0_Im : mem_17_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_18 = 5'h12 == io_in_waddr_0 ? io_in_data_0_Im : mem_18_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_19 = 5'h13 == io_in_waddr_0 ? io_in_data_0_Im : mem_19_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_20 = 5'h14 == io_in_waddr_0 ? io_in_data_0_Im : mem_20_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_21 = 5'h15 == io_in_waddr_0 ? io_in_data_0_Im : mem_21_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_22 = 5'h16 == io_in_waddr_0 ? io_in_data_0_Im : mem_22_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_23 = 5'h17 == io_in_waddr_0 ? io_in_data_0_Im : mem_23_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_24 = 5'h0 == io_in_waddr_0 ? io_in_data_0_Re : mem_0_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_25 = 5'h1 == io_in_waddr_0 ? io_in_data_0_Re : mem_1_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_26 = 5'h2 == io_in_waddr_0 ? io_in_data_0_Re : mem_2_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_27 = 5'h3 == io_in_waddr_0 ? io_in_data_0_Re : mem_3_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_28 = 5'h4 == io_in_waddr_0 ? io_in_data_0_Re : mem_4_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_29 = 5'h5 == io_in_waddr_0 ? io_in_data_0_Re : mem_5_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_30 = 5'h6 == io_in_waddr_0 ? io_in_data_0_Re : mem_6_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_31 = 5'h7 == io_in_waddr_0 ? io_in_data_0_Re : mem_7_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_32 = 5'h8 == io_in_waddr_0 ? io_in_data_0_Re : mem_8_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_33 = 5'h9 == io_in_waddr_0 ? io_in_data_0_Re : mem_9_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_34 = 5'ha == io_in_waddr_0 ? io_in_data_0_Re : mem_10_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_35 = 5'hb == io_in_waddr_0 ? io_in_data_0_Re : mem_11_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_36 = 5'hc == io_in_waddr_0 ? io_in_data_0_Re : mem_12_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_37 = 5'hd == io_in_waddr_0 ? io_in_data_0_Re : mem_13_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_38 = 5'he == io_in_waddr_0 ? io_in_data_0_Re : mem_14_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_39 = 5'hf == io_in_waddr_0 ? io_in_data_0_Re : mem_15_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_40 = 5'h10 == io_in_waddr_0 ? io_in_data_0_Re : mem_16_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_41 = 5'h11 == io_in_waddr_0 ? io_in_data_0_Re : mem_17_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_42 = 5'h12 == io_in_waddr_0 ? io_in_data_0_Re : mem_18_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_43 = 5'h13 == io_in_waddr_0 ? io_in_data_0_Re : mem_19_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_44 = 5'h14 == io_in_waddr_0 ? io_in_data_0_Re : mem_20_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_45 = 5'h15 == io_in_waddr_0 ? io_in_data_0_Re : mem_21_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_46 = 5'h16 == io_in_waddr_0 ? io_in_data_0_Re : mem_22_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_47 = 5'h17 == io_in_waddr_0 ? io_in_data_0_Re : mem_23_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_48 = io_wr_0 ? _GEN_0 : mem_0_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_49 = io_wr_0 ? _GEN_1 : mem_1_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_50 = io_wr_0 ? _GEN_2 : mem_2_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_51 = io_wr_0 ? _GEN_3 : mem_3_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_52 = io_wr_0 ? _GEN_4 : mem_4_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_53 = io_wr_0 ? _GEN_5 : mem_5_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_54 = io_wr_0 ? _GEN_6 : mem_6_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_55 = io_wr_0 ? _GEN_7 : mem_7_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_56 = io_wr_0 ? _GEN_8 : mem_8_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_57 = io_wr_0 ? _GEN_9 : mem_9_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_58 = io_wr_0 ? _GEN_10 : mem_10_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_59 = io_wr_0 ? _GEN_11 : mem_11_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_60 = io_wr_0 ? _GEN_12 : mem_12_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_61 = io_wr_0 ? _GEN_13 : mem_13_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_62 = io_wr_0 ? _GEN_14 : mem_14_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_63 = io_wr_0 ? _GEN_15 : mem_15_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_64 = io_wr_0 ? _GEN_16 : mem_16_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_65 = io_wr_0 ? _GEN_17 : mem_17_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_66 = io_wr_0 ? _GEN_18 : mem_18_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_67 = io_wr_0 ? _GEN_19 : mem_19_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_68 = io_wr_0 ? _GEN_20 : mem_20_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_69 = io_wr_0 ? _GEN_21 : mem_21_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_70 = io_wr_0 ? _GEN_22 : mem_22_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_71 = io_wr_0 ? _GEN_23 : mem_23_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_72 = io_wr_0 ? _GEN_24 : mem_0_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_73 = io_wr_0 ? _GEN_25 : mem_1_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_74 = io_wr_0 ? _GEN_26 : mem_2_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_75 = io_wr_0 ? _GEN_27 : mem_3_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_76 = io_wr_0 ? _GEN_28 : mem_4_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_77 = io_wr_0 ? _GEN_29 : mem_5_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_78 = io_wr_0 ? _GEN_30 : mem_6_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_79 = io_wr_0 ? _GEN_31 : mem_7_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_80 = io_wr_0 ? _GEN_32 : mem_8_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_81 = io_wr_0 ? _GEN_33 : mem_9_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_82 = io_wr_0 ? _GEN_34 : mem_10_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_83 = io_wr_0 ? _GEN_35 : mem_11_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_84 = io_wr_0 ? _GEN_36 : mem_12_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_85 = io_wr_0 ? _GEN_37 : mem_13_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_86 = io_wr_0 ? _GEN_38 : mem_14_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_87 = io_wr_0 ? _GEN_39 : mem_15_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_88 = io_wr_0 ? _GEN_40 : mem_16_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_89 = io_wr_0 ? _GEN_41 : mem_17_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_90 = io_wr_0 ? _GEN_42 : mem_18_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_91 = io_wr_0 ? _GEN_43 : mem_19_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_92 = io_wr_0 ? _GEN_44 : mem_20_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_93 = io_wr_0 ? _GEN_45 : mem_21_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_94 = io_wr_0 ? _GEN_46 : mem_22_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_95 = io_wr_0 ? _GEN_47 : mem_23_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_193 = 5'h1 == io_in_raddr ? mem_1_Im : mem_0_Im; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_194 = 5'h2 == io_in_raddr ? mem_2_Im : _GEN_193; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_195 = 5'h3 == io_in_raddr ? mem_3_Im : _GEN_194; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_196 = 5'h4 == io_in_raddr ? mem_4_Im : _GEN_195; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_197 = 5'h5 == io_in_raddr ? mem_5_Im : _GEN_196; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_198 = 5'h6 == io_in_raddr ? mem_6_Im : _GEN_197; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_199 = 5'h7 == io_in_raddr ? mem_7_Im : _GEN_198; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_200 = 5'h8 == io_in_raddr ? mem_8_Im : _GEN_199; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_201 = 5'h9 == io_in_raddr ? mem_9_Im : _GEN_200; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_202 = 5'ha == io_in_raddr ? mem_10_Im : _GEN_201; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_203 = 5'hb == io_in_raddr ? mem_11_Im : _GEN_202; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_204 = 5'hc == io_in_raddr ? mem_12_Im : _GEN_203; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_205 = 5'hd == io_in_raddr ? mem_13_Im : _GEN_204; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_206 = 5'he == io_in_raddr ? mem_14_Im : _GEN_205; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_207 = 5'hf == io_in_raddr ? mem_15_Im : _GEN_206; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_208 = 5'h10 == io_in_raddr ? mem_16_Im : _GEN_207; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_209 = 5'h11 == io_in_raddr ? mem_17_Im : _GEN_208; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_210 = 5'h12 == io_in_raddr ? mem_18_Im : _GEN_209; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_211 = 5'h13 == io_in_raddr ? mem_19_Im : _GEN_210; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_212 = 5'h14 == io_in_raddr ? mem_20_Im : _GEN_211; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_213 = 5'h15 == io_in_raddr ? mem_21_Im : _GEN_212; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_214 = 5'h16 == io_in_raddr ? mem_22_Im : _GEN_213; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_215 = 5'h17 == io_in_raddr ? mem_23_Im : _GEN_214; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_217 = 5'h1 == io_in_raddr ? mem_1_Re : mem_0_Re; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_218 = 5'h2 == io_in_raddr ? mem_2_Re : _GEN_217; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_219 = 5'h3 == io_in_raddr ? mem_3_Re : _GEN_218; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_220 = 5'h4 == io_in_raddr ? mem_4_Re : _GEN_219; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_221 = 5'h5 == io_in_raddr ? mem_5_Re : _GEN_220; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_222 = 5'h6 == io_in_raddr ? mem_6_Re : _GEN_221; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_223 = 5'h7 == io_in_raddr ? mem_7_Re : _GEN_222; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_224 = 5'h8 == io_in_raddr ? mem_8_Re : _GEN_223; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_225 = 5'h9 == io_in_raddr ? mem_9_Re : _GEN_224; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_226 = 5'ha == io_in_raddr ? mem_10_Re : _GEN_225; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_227 = 5'hb == io_in_raddr ? mem_11_Re : _GEN_226; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_228 = 5'hc == io_in_raddr ? mem_12_Re : _GEN_227; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_229 = 5'hd == io_in_raddr ? mem_13_Re : _GEN_228; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_230 = 5'he == io_in_raddr ? mem_14_Re : _GEN_229; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_231 = 5'hf == io_in_raddr ? mem_15_Re : _GEN_230; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_232 = 5'h10 == io_in_raddr ? mem_16_Re : _GEN_231; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_233 = 5'h11 == io_in_raddr ? mem_17_Re : _GEN_232; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_234 = 5'h12 == io_in_raddr ? mem_18_Re : _GEN_233; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_235 = 5'h13 == io_in_raddr ? mem_19_Re : _GEN_234; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_236 = 5'h14 == io_in_raddr ? mem_20_Re : _GEN_235; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_237 = 5'h15 == io_in_raddr ? mem_21_Re : _GEN_236; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_238 = 5'h16 == io_in_raddr ? mem_22_Re : _GEN_237; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_239 = 5'h17 == io_in_raddr ? mem_23_Re : _GEN_238; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_240 = io_re ? _GEN_215 : 32'h0; // @[FFTDesigns.scala 3320:18 3321:21 3324:24]
  wire [31:0] _GEN_241 = io_re ? _GEN_239 : 32'h0; // @[FFTDesigns.scala 3320:18 3321:21 3323:24]
  assign io_out_data_Re = io_en ? _GEN_241 : 32'h0; // @[FFTDesigns.scala 3314:16 3327:22]
  assign io_out_data_Im = io_en ? _GEN_240 : 32'h0; // @[FFTDesigns.scala 3314:16 3328:22]
  always @(posedge clock) begin
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h0 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_0_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_0_Re <= _GEN_72;
        end
      end else begin
        mem_0_Re <= _GEN_72;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h0 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_0_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_0_Im <= _GEN_48;
        end
      end else begin
        mem_0_Im <= _GEN_48;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h1 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_1_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_1_Re <= _GEN_73;
        end
      end else begin
        mem_1_Re <= _GEN_73;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h1 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_1_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_1_Im <= _GEN_49;
        end
      end else begin
        mem_1_Im <= _GEN_49;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h2 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_2_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_2_Re <= _GEN_74;
        end
      end else begin
        mem_2_Re <= _GEN_74;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h2 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_2_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_2_Im <= _GEN_50;
        end
      end else begin
        mem_2_Im <= _GEN_50;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h3 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_3_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_3_Re <= _GEN_75;
        end
      end else begin
        mem_3_Re <= _GEN_75;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h3 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_3_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_3_Im <= _GEN_51;
        end
      end else begin
        mem_3_Im <= _GEN_51;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h4 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_4_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_4_Re <= _GEN_76;
        end
      end else begin
        mem_4_Re <= _GEN_76;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h4 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_4_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_4_Im <= _GEN_52;
        end
      end else begin
        mem_4_Im <= _GEN_52;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h5 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_5_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_5_Re <= _GEN_77;
        end
      end else begin
        mem_5_Re <= _GEN_77;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h5 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_5_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_5_Im <= _GEN_53;
        end
      end else begin
        mem_5_Im <= _GEN_53;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h6 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_6_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_6_Re <= _GEN_78;
        end
      end else begin
        mem_6_Re <= _GEN_78;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h6 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_6_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_6_Im <= _GEN_54;
        end
      end else begin
        mem_6_Im <= _GEN_54;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h7 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_7_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_7_Re <= _GEN_79;
        end
      end else begin
        mem_7_Re <= _GEN_79;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h7 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_7_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_7_Im <= _GEN_55;
        end
      end else begin
        mem_7_Im <= _GEN_55;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h8 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_8_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_8_Re <= _GEN_80;
        end
      end else begin
        mem_8_Re <= _GEN_80;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h8 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_8_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_8_Im <= _GEN_56;
        end
      end else begin
        mem_8_Im <= _GEN_56;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h9 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_9_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_9_Re <= _GEN_81;
        end
      end else begin
        mem_9_Re <= _GEN_81;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h9 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_9_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_9_Im <= _GEN_57;
        end
      end else begin
        mem_9_Im <= _GEN_57;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'ha == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_10_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_10_Re <= _GEN_82;
        end
      end else begin
        mem_10_Re <= _GEN_82;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'ha == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_10_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_10_Im <= _GEN_58;
        end
      end else begin
        mem_10_Im <= _GEN_58;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'hb == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_11_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_11_Re <= _GEN_83;
        end
      end else begin
        mem_11_Re <= _GEN_83;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'hb == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_11_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_11_Im <= _GEN_59;
        end
      end else begin
        mem_11_Im <= _GEN_59;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'hc == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_12_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_12_Re <= _GEN_84;
        end
      end else begin
        mem_12_Re <= _GEN_84;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'hc == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_12_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_12_Im <= _GEN_60;
        end
      end else begin
        mem_12_Im <= _GEN_60;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'hd == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_13_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_13_Re <= _GEN_85;
        end
      end else begin
        mem_13_Re <= _GEN_85;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'hd == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_13_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_13_Im <= _GEN_61;
        end
      end else begin
        mem_13_Im <= _GEN_61;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'he == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_14_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_14_Re <= _GEN_86;
        end
      end else begin
        mem_14_Re <= _GEN_86;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'he == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_14_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_14_Im <= _GEN_62;
        end
      end else begin
        mem_14_Im <= _GEN_62;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'hf == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_15_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_15_Re <= _GEN_87;
        end
      end else begin
        mem_15_Re <= _GEN_87;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'hf == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_15_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_15_Im <= _GEN_63;
        end
      end else begin
        mem_15_Im <= _GEN_63;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h10 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_16_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_16_Re <= _GEN_88;
        end
      end else begin
        mem_16_Re <= _GEN_88;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h10 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_16_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_16_Im <= _GEN_64;
        end
      end else begin
        mem_16_Im <= _GEN_64;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h11 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_17_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_17_Re <= _GEN_89;
        end
      end else begin
        mem_17_Re <= _GEN_89;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h11 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_17_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_17_Im <= _GEN_65;
        end
      end else begin
        mem_17_Im <= _GEN_65;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h12 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_18_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_18_Re <= _GEN_90;
        end
      end else begin
        mem_18_Re <= _GEN_90;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h12 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_18_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_18_Im <= _GEN_66;
        end
      end else begin
        mem_18_Im <= _GEN_66;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h13 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_19_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_19_Re <= _GEN_91;
        end
      end else begin
        mem_19_Re <= _GEN_91;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h13 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_19_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_19_Im <= _GEN_67;
        end
      end else begin
        mem_19_Im <= _GEN_67;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h14 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_20_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_20_Re <= _GEN_92;
        end
      end else begin
        mem_20_Re <= _GEN_92;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h14 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_20_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_20_Im <= _GEN_68;
        end
      end else begin
        mem_20_Im <= _GEN_68;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h15 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_21_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_21_Re <= _GEN_93;
        end
      end else begin
        mem_21_Re <= _GEN_93;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h15 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_21_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_21_Im <= _GEN_69;
        end
      end else begin
        mem_21_Im <= _GEN_69;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h16 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_22_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_22_Re <= _GEN_94;
        end
      end else begin
        mem_22_Re <= _GEN_94;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h16 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_22_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_22_Im <= _GEN_70;
        end
      end else begin
        mem_22_Im <= _GEN_70;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h17 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_23_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_23_Re <= _GEN_95;
        end
      end else begin
        mem_23_Re <= _GEN_95;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (5'h17 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_23_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_23_Im <= _GEN_71;
        end
      end else begin
        mem_23_Im <= _GEN_71;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_3_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_4_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_4_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_5_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_5_Im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_6_Re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_6_Im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_7_Re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_7_Im = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mem_8_Re = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mem_8_Im = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_9_Re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mem_9_Im = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mem_10_Re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mem_10_Im = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_11_Re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mem_11_Im = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  mem_12_Re = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  mem_12_Im = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  mem_13_Re = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mem_13_Im = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mem_14_Re = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  mem_14_Im = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  mem_15_Re = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  mem_15_Im = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mem_16_Re = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mem_16_Im = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mem_17_Re = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  mem_17_Im = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  mem_18_Re = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  mem_18_Im = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  mem_19_Re = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  mem_19_Im = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  mem_20_Re = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  mem_20_Im = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  mem_21_Re = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  mem_21_Im = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  mem_22_Re = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  mem_22_Im = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  mem_23_Re = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  mem_23_Im = _RAND_47[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PermutationsWithStreaming_mr_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  input         io_in_en_5,
  input         io_in_en_6,
  input         io_in_en_7,
  input         io_in_en_8,
  input         io_in_en_9,
  input         io_in_en_10,
  input         io_in_en_11,
  input         io_in_en_12,
  input         io_in_en_13,
  input         io_in_en_14,
  input         io_in_en_15,
  input         io_in_en_16,
  input         io_in_en_17,
  input         io_in_en_18,
  input         io_in_en_19,
  input         io_in_en_20,
  input         io_in_en_21,
  input         io_in_en_22,
  input         io_in_en_23,
  input         io_in_en_24,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_mw_clock; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_clock; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_1_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_1_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_1_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_clock; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_2_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_2_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_2_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_clock; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_3_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_3_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_3_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_clock; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_4_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_4_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_4_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_clock; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_5_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_5_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_5_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_clock; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_6_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_6_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_6_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_clock; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_7_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_7_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [4:0] RAM_Block_mw_7_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [4:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2907:28]
  wire [2:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2907:28]
  wire [2:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2907:28]
  wire [2:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2907:28]
  wire [2:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2907:28]
  wire [2:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2907:28]
  wire [2:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2907:28]
  wire [2:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2907:28]
  wire [3:0] M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2908:29]
  wire [4:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2908:29]
  wire [4:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2908:29]
  wire [4:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2908:29]
  wire [4:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2908:29]
  wire [4:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2908:29]
  wire [4:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2908:29]
  wire [4:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2908:29]
  wire [4:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2909:29]
  wire [4:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2909:29]
  wire [4:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2909:29]
  wire [4:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2909:29]
  wire [4:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2909:29]
  wire [4:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2909:29]
  wire [4:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2909:29]
  wire [4:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2909:29]
  wire [4:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2909:29]
  wire [3:0] Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2910:31]
  wire [2:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2910:31]
  wire [2:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2910:31]
  wire [2:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2910:31]
  wire [2:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2910:31]
  wire [2:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2910:31]
  wire [2:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2910:31]
  wire [2:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2910:31]
  reg  offset_switch; // @[FFTDesigns.scala 2710:28]
  reg [31:0] input_delay_registers_0_0_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_0_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_1_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_1_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_2_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_2_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_3_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_3_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_4_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_4_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_5_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_5_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_6_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_6_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_7_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_7_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_8_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_8_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_9_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_9_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_10_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_10_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_11_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_11_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_1_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_1_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_2_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_2_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_3_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_3_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_4_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_4_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_5_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_5_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_6_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_6_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_7_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_7_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_8_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_8_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_9_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_9_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_10_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_10_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_11_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_11_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_0_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_0_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_1_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_1_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_2_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_2_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_3_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_3_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_4_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_4_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_5_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_5_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_6_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_6_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_7_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_7_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_8_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_8_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_9_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_9_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_10_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_10_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_11_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_2_11_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_1_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_1_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_2_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_2_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_3_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_3_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_4_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_4_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_5_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_5_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_6_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_6_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_7_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_7_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_8_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_8_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_9_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_9_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_10_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_10_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_11_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_3_11_Im; // @[FFTDesigns.scala 2834:42]
  reg [3:0] cnt2; // @[FFTDesigns.scala 2912:25]
  reg [2:0] cnt; // @[FFTDesigns.scala 2913:24]
  wire [5:0] lo_lo = {io_in_en_5,io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2914:21]
  wire [11:0] lo = {io_in_en_11,io_in_en_10,io_in_en_9,io_in_en_8,io_in_en_7,io_in_en_6,lo_lo}; // @[FFTDesigns.scala 2914:21]
  wire [5:0] hi_lo = {io_in_en_17,io_in_en_16,io_in_en_15,io_in_en_14,io_in_en_13,io_in_en_12}; // @[FFTDesigns.scala 2914:21]
  wire [24:0] _T = {io_in_en_24,io_in_en_23,io_in_en_22,io_in_en_21,io_in_en_20,io_in_en_19,io_in_en_18,hi_lo,lo}; // @[FFTDesigns.scala 2914:21]
  wire  M0_0_re = |_T; // @[FFTDesigns.scala 2914:28]
  wire  _T_3 = cnt == 3'h7; // @[FFTDesigns.scala 2922:46]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2925:28]
  wire [3:0] _cnt2_T_1 = cnt2 + 4'h1; // @[FFTDesigns.scala 2928:24]
  wire [2:0] _cnt_T_1 = cnt + 3'h1; // @[FFTDesigns.scala 2933:24]
  wire [2:0] _GEN_0 = cnt2 >= 4'h4 ? _cnt_T_1 : 3'h0; // @[FFTDesigns.scala 2932:32 2933:17 2935:17]
  wire  _GEN_6 = cnt2 == 4'hb & cnt == 3'h7 ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2922:69 2925:25]
  wire [4:0] _M0_0_in_raddr_T_1 = 4'hc * _offset_switch_T; // @[FFTDesigns.scala 2950:56]
  wire [4:0] _M0_0_in_raddr_T_3 = M0_Config_ROM_io_out_0 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [4:0] _GEN_1024 = {{1'd0}, cnt2}; // @[FFTDesigns.scala 2951:34]
  wire [4:0] _M1_0_in_raddr_T_3 = _GEN_1024 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2951:34]
  wire [4:0] _M1_0_in_waddr_T = 4'hc * offset_switch; // @[FFTDesigns.scala 2952:56]
  wire [4:0] _M1_0_in_waddr_T_2 = M1_Config_ROM_io_out_0 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [4:0] _M0_1_in_raddr_T_3 = M0_Config_ROM_io_out_1 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [4:0] _M1_1_in_waddr_T_2 = M1_Config_ROM_io_out_1 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [4:0] _M0_2_in_raddr_T_3 = M0_Config_ROM_io_out_2 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [4:0] _M1_2_in_waddr_T_2 = M1_Config_ROM_io_out_2 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [4:0] _M0_3_in_raddr_T_3 = M0_Config_ROM_io_out_3 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [4:0] _M1_3_in_waddr_T_2 = M1_Config_ROM_io_out_3 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [4:0] _M0_4_in_raddr_T_3 = M0_Config_ROM_io_out_4 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [4:0] _M1_4_in_waddr_T_2 = M1_Config_ROM_io_out_4 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [4:0] _M0_5_in_raddr_T_3 = M0_Config_ROM_io_out_5 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [4:0] _M1_5_in_waddr_T_2 = M1_Config_ROM_io_out_5 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [4:0] _M0_6_in_raddr_T_3 = M0_Config_ROM_io_out_6 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [4:0] _M1_6_in_waddr_T_2 = M1_Config_ROM_io_out_6 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [4:0] _M0_7_in_raddr_T_3 = M0_Config_ROM_io_out_7 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [4:0] _M1_7_in_waddr_T_2 = M1_Config_ROM_io_out_7 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _GEN_16 = 3'h1 == cnt ? 4'h2 : 4'h0; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_17 = 3'h2 == cnt ? 4'h3 : _GEN_16; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_18 = 3'h3 == cnt ? 4'h5 : _GEN_17; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_19 = 3'h4 == cnt ? 4'h6 : _GEN_18; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_20 = 3'h5 == cnt ? 4'h8 : _GEN_19; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_21 = 3'h6 == cnt ? 4'h9 : _GEN_20; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_22 = 3'h7 == cnt ? 4'hb : _GEN_21; // @[FFTDesigns.scala 2978:{55,55}]
  wire [4:0] _GEN_1032 = {{1'd0}, _GEN_22}; // @[FFTDesigns.scala 2978:55]
  wire [4:0] _M0_0_in_waddr_0_T_2 = _GEN_1032 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2978:55]
  wire [3:0] _GEN_24 = 3'h1 == cnt ? 4'h4 : 4'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_25 = 3'h2 == cnt ? 4'h0 : _GEN_24; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_26 = 3'h3 == cnt ? 4'h4 : _GEN_25; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_27 = 3'h4 == cnt ? 4'h0 : _GEN_26; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_28 = 3'h5 == cnt ? 4'h4 : _GEN_27; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_29 = 3'h6 == cnt ? 4'h0 : _GEN_28; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_30 = 3'h7 == cnt ? 4'h4 : _GEN_29; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_32 = 4'h1 == _GEN_30 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_33 = 4'h2 == _GEN_30 ? input_delay_registers_3_2_Im : _GEN_32; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_34 = 4'h3 == _GEN_30 ? input_delay_registers_3_3_Im : _GEN_33; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_35 = 4'h4 == _GEN_30 ? input_delay_registers_3_4_Im : _GEN_34; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_36 = 4'h5 == _GEN_30 ? input_delay_registers_3_5_Im : _GEN_35; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_37 = 4'h6 == _GEN_30 ? input_delay_registers_3_6_Im : _GEN_36; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_38 = 4'h7 == _GEN_30 ? input_delay_registers_3_7_Im : _GEN_37; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_39 = 4'h8 == _GEN_30 ? input_delay_registers_3_8_Im : _GEN_38; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_40 = 4'h9 == _GEN_30 ? input_delay_registers_3_9_Im : _GEN_39; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_41 = 4'ha == _GEN_30 ? input_delay_registers_3_10_Im : _GEN_40; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_42 = 4'hb == _GEN_30 ? input_delay_registers_3_11_Im : _GEN_41; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_44 = 4'h1 == _GEN_30 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_45 = 4'h2 == _GEN_30 ? input_delay_registers_3_2_Re : _GEN_44; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_46 = 4'h3 == _GEN_30 ? input_delay_registers_3_3_Re : _GEN_45; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_47 = 4'h4 == _GEN_30 ? input_delay_registers_3_4_Re : _GEN_46; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_48 = 4'h5 == _GEN_30 ? input_delay_registers_3_5_Re : _GEN_47; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_49 = 4'h6 == _GEN_30 ? input_delay_registers_3_6_Re : _GEN_48; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_50 = 4'h7 == _GEN_30 ? input_delay_registers_3_7_Re : _GEN_49; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_51 = 4'h8 == _GEN_30 ? input_delay_registers_3_8_Re : _GEN_50; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_52 = 4'h9 == _GEN_30 ? input_delay_registers_3_9_Re : _GEN_51; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_53 = 4'ha == _GEN_30 ? input_delay_registers_3_10_Re : _GEN_52; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_54 = 4'hb == _GEN_30 ? input_delay_registers_3_11_Re : _GEN_53; // @[FFTDesigns.scala 2979:{32,32}]
  wire  _GEN_56 = 3'h1 == cnt ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2977:{27,27}]
  wire  _GEN_58 = 3'h3 == cnt ? 1'h0 : 3'h2 == cnt | _GEN_56; // @[FFTDesigns.scala 2977:{27,27}]
  wire  _GEN_60 = 3'h5 == cnt ? 1'h0 : 3'h4 == cnt | _GEN_58; // @[FFTDesigns.scala 2977:{27,27}]
  wire  _GEN_62 = 3'h7 == cnt ? 1'h0 : 3'h6 == cnt | _GEN_60; // @[FFTDesigns.scala 2977:{27,27}]
  wire [3:0] _GEN_64 = 3'h1 == cnt ? 4'h0 : 4'h1; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_65 = 3'h2 == cnt ? 4'h4 : _GEN_64; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_66 = 3'h3 == cnt ? 4'h0 : _GEN_65; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_67 = 3'h4 == cnt ? 4'h7 : _GEN_66; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_68 = 3'h5 == cnt ? 4'h0 : _GEN_67; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_69 = 3'h6 == cnt ? 4'ha : _GEN_68; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_70 = 3'h7 == cnt ? 4'h0 : _GEN_69; // @[FFTDesigns.scala 2978:{55,55}]
  wire [4:0] _GEN_1036 = {{1'd0}, _GEN_70}; // @[FFTDesigns.scala 2978:55]
  wire [4:0] _M0_0_in_waddr_1_T_2 = _GEN_1036 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2978:55]
  wire [3:0] _GEN_72 = 3'h1 == cnt ? 4'h0 : 4'h8; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_73 = 3'h2 == cnt ? 4'h8 : _GEN_72; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_74 = 3'h3 == cnt ? 4'h0 : _GEN_73; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_75 = 3'h4 == cnt ? 4'h8 : _GEN_74; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_76 = 3'h5 == cnt ? 4'h0 : _GEN_75; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_77 = 3'h6 == cnt ? 4'h8 : _GEN_76; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_78 = 3'h7 == cnt ? 4'h0 : _GEN_77; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_80 = 4'h1 == _GEN_78 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_81 = 4'h2 == _GEN_78 ? input_delay_registers_3_2_Im : _GEN_80; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_82 = 4'h3 == _GEN_78 ? input_delay_registers_3_3_Im : _GEN_81; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_83 = 4'h4 == _GEN_78 ? input_delay_registers_3_4_Im : _GEN_82; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_84 = 4'h5 == _GEN_78 ? input_delay_registers_3_5_Im : _GEN_83; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_85 = 4'h6 == _GEN_78 ? input_delay_registers_3_6_Im : _GEN_84; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_86 = 4'h7 == _GEN_78 ? input_delay_registers_3_7_Im : _GEN_85; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_87 = 4'h8 == _GEN_78 ? input_delay_registers_3_8_Im : _GEN_86; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_88 = 4'h9 == _GEN_78 ? input_delay_registers_3_9_Im : _GEN_87; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_89 = 4'ha == _GEN_78 ? input_delay_registers_3_10_Im : _GEN_88; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_90 = 4'hb == _GEN_78 ? input_delay_registers_3_11_Im : _GEN_89; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_92 = 4'h1 == _GEN_78 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_93 = 4'h2 == _GEN_78 ? input_delay_registers_3_2_Re : _GEN_92; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_94 = 4'h3 == _GEN_78 ? input_delay_registers_3_3_Re : _GEN_93; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_95 = 4'h4 == _GEN_78 ? input_delay_registers_3_4_Re : _GEN_94; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_96 = 4'h5 == _GEN_78 ? input_delay_registers_3_5_Re : _GEN_95; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_97 = 4'h6 == _GEN_78 ? input_delay_registers_3_6_Re : _GEN_96; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_98 = 4'h7 == _GEN_78 ? input_delay_registers_3_7_Re : _GEN_97; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_99 = 4'h8 == _GEN_78 ? input_delay_registers_3_8_Re : _GEN_98; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_100 = 4'h9 == _GEN_78 ? input_delay_registers_3_9_Re : _GEN_99; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_101 = 4'ha == _GEN_78 ? input_delay_registers_3_10_Re : _GEN_100; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_102 = 4'hb == _GEN_78 ? input_delay_registers_3_11_Re : _GEN_101; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_120 = 3'h1 == cnt ? 4'h5 : 4'h1; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_121 = 3'h2 == cnt ? 4'h1 : _GEN_120; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_122 = 3'h3 == cnt ? 4'h5 : _GEN_121; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_123 = 3'h4 == cnt ? 4'h1 : _GEN_122; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_124 = 3'h5 == cnt ? 4'h5 : _GEN_123; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_125 = 3'h6 == cnt ? 4'h1 : _GEN_124; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_126 = 3'h7 == cnt ? 4'h5 : _GEN_125; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_128 = 4'h1 == _GEN_126 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_129 = 4'h2 == _GEN_126 ? input_delay_registers_3_2_Im : _GEN_128; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_130 = 4'h3 == _GEN_126 ? input_delay_registers_3_3_Im : _GEN_129; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_131 = 4'h4 == _GEN_126 ? input_delay_registers_3_4_Im : _GEN_130; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_132 = 4'h5 == _GEN_126 ? input_delay_registers_3_5_Im : _GEN_131; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_133 = 4'h6 == _GEN_126 ? input_delay_registers_3_6_Im : _GEN_132; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_134 = 4'h7 == _GEN_126 ? input_delay_registers_3_7_Im : _GEN_133; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_135 = 4'h8 == _GEN_126 ? input_delay_registers_3_8_Im : _GEN_134; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_136 = 4'h9 == _GEN_126 ? input_delay_registers_3_9_Im : _GEN_135; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_137 = 4'ha == _GEN_126 ? input_delay_registers_3_10_Im : _GEN_136; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_138 = 4'hb == _GEN_126 ? input_delay_registers_3_11_Im : _GEN_137; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_140 = 4'h1 == _GEN_126 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_141 = 4'h2 == _GEN_126 ? input_delay_registers_3_2_Re : _GEN_140; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_142 = 4'h3 == _GEN_126 ? input_delay_registers_3_3_Re : _GEN_141; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_143 = 4'h4 == _GEN_126 ? input_delay_registers_3_4_Re : _GEN_142; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_144 = 4'h5 == _GEN_126 ? input_delay_registers_3_5_Re : _GEN_143; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_145 = 4'h6 == _GEN_126 ? input_delay_registers_3_6_Re : _GEN_144; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_146 = 4'h7 == _GEN_126 ? input_delay_registers_3_7_Re : _GEN_145; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_147 = 4'h8 == _GEN_126 ? input_delay_registers_3_8_Re : _GEN_146; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_148 = 4'h9 == _GEN_126 ? input_delay_registers_3_9_Re : _GEN_147; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_149 = 4'ha == _GEN_126 ? input_delay_registers_3_10_Re : _GEN_148; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_150 = 4'hb == _GEN_126 ? input_delay_registers_3_11_Re : _GEN_149; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_168 = 3'h1 == cnt ? 4'h0 : 4'h9; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_169 = 3'h2 == cnt ? 4'h9 : _GEN_168; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_170 = 3'h3 == cnt ? 4'h0 : _GEN_169; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_171 = 3'h4 == cnt ? 4'h9 : _GEN_170; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_172 = 3'h5 == cnt ? 4'h0 : _GEN_171; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_173 = 3'h6 == cnt ? 4'h9 : _GEN_172; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_174 = 3'h7 == cnt ? 4'h0 : _GEN_173; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_176 = 4'h1 == _GEN_174 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_177 = 4'h2 == _GEN_174 ? input_delay_registers_3_2_Im : _GEN_176; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_178 = 4'h3 == _GEN_174 ? input_delay_registers_3_3_Im : _GEN_177; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_179 = 4'h4 == _GEN_174 ? input_delay_registers_3_4_Im : _GEN_178; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_180 = 4'h5 == _GEN_174 ? input_delay_registers_3_5_Im : _GEN_179; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_181 = 4'h6 == _GEN_174 ? input_delay_registers_3_6_Im : _GEN_180; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_182 = 4'h7 == _GEN_174 ? input_delay_registers_3_7_Im : _GEN_181; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_183 = 4'h8 == _GEN_174 ? input_delay_registers_3_8_Im : _GEN_182; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_184 = 4'h9 == _GEN_174 ? input_delay_registers_3_9_Im : _GEN_183; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_185 = 4'ha == _GEN_174 ? input_delay_registers_3_10_Im : _GEN_184; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_186 = 4'hb == _GEN_174 ? input_delay_registers_3_11_Im : _GEN_185; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_188 = 4'h1 == _GEN_174 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_189 = 4'h2 == _GEN_174 ? input_delay_registers_3_2_Re : _GEN_188; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_190 = 4'h3 == _GEN_174 ? input_delay_registers_3_3_Re : _GEN_189; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_191 = 4'h4 == _GEN_174 ? input_delay_registers_3_4_Re : _GEN_190; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_192 = 4'h5 == _GEN_174 ? input_delay_registers_3_5_Re : _GEN_191; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_193 = 4'h6 == _GEN_174 ? input_delay_registers_3_6_Re : _GEN_192; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_194 = 4'h7 == _GEN_174 ? input_delay_registers_3_7_Re : _GEN_193; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_195 = 4'h8 == _GEN_174 ? input_delay_registers_3_8_Re : _GEN_194; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_196 = 4'h9 == _GEN_174 ? input_delay_registers_3_9_Re : _GEN_195; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_197 = 4'ha == _GEN_174 ? input_delay_registers_3_10_Re : _GEN_196; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_198 = 4'hb == _GEN_174 ? input_delay_registers_3_11_Re : _GEN_197; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_216 = 3'h1 == cnt ? 4'h6 : 4'h2; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_217 = 3'h2 == cnt ? 4'h2 : _GEN_216; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_218 = 3'h3 == cnt ? 4'h6 : _GEN_217; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_219 = 3'h4 == cnt ? 4'h2 : _GEN_218; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_220 = 3'h5 == cnt ? 4'h6 : _GEN_219; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_221 = 3'h6 == cnt ? 4'h2 : _GEN_220; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_222 = 3'h7 == cnt ? 4'h6 : _GEN_221; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_224 = 4'h1 == _GEN_222 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_225 = 4'h2 == _GEN_222 ? input_delay_registers_3_2_Im : _GEN_224; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_226 = 4'h3 == _GEN_222 ? input_delay_registers_3_3_Im : _GEN_225; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_227 = 4'h4 == _GEN_222 ? input_delay_registers_3_4_Im : _GEN_226; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_228 = 4'h5 == _GEN_222 ? input_delay_registers_3_5_Im : _GEN_227; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_229 = 4'h6 == _GEN_222 ? input_delay_registers_3_6_Im : _GEN_228; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_230 = 4'h7 == _GEN_222 ? input_delay_registers_3_7_Im : _GEN_229; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_231 = 4'h8 == _GEN_222 ? input_delay_registers_3_8_Im : _GEN_230; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_232 = 4'h9 == _GEN_222 ? input_delay_registers_3_9_Im : _GEN_231; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_233 = 4'ha == _GEN_222 ? input_delay_registers_3_10_Im : _GEN_232; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_234 = 4'hb == _GEN_222 ? input_delay_registers_3_11_Im : _GEN_233; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_236 = 4'h1 == _GEN_222 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_237 = 4'h2 == _GEN_222 ? input_delay_registers_3_2_Re : _GEN_236; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_238 = 4'h3 == _GEN_222 ? input_delay_registers_3_3_Re : _GEN_237; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_239 = 4'h4 == _GEN_222 ? input_delay_registers_3_4_Re : _GEN_238; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_240 = 4'h5 == _GEN_222 ? input_delay_registers_3_5_Re : _GEN_239; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_241 = 4'h6 == _GEN_222 ? input_delay_registers_3_6_Re : _GEN_240; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_242 = 4'h7 == _GEN_222 ? input_delay_registers_3_7_Re : _GEN_241; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_243 = 4'h8 == _GEN_222 ? input_delay_registers_3_8_Re : _GEN_242; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_244 = 4'h9 == _GEN_222 ? input_delay_registers_3_9_Re : _GEN_243; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_245 = 4'ha == _GEN_222 ? input_delay_registers_3_10_Re : _GEN_244; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_246 = 4'hb == _GEN_222 ? input_delay_registers_3_11_Re : _GEN_245; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_264 = 3'h1 == cnt ? 4'h0 : 4'ha; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_265 = 3'h2 == cnt ? 4'ha : _GEN_264; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_266 = 3'h3 == cnt ? 4'h0 : _GEN_265; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_267 = 3'h4 == cnt ? 4'ha : _GEN_266; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_268 = 3'h5 == cnt ? 4'h0 : _GEN_267; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_269 = 3'h6 == cnt ? 4'ha : _GEN_268; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_270 = 3'h7 == cnt ? 4'h0 : _GEN_269; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_272 = 4'h1 == _GEN_270 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_273 = 4'h2 == _GEN_270 ? input_delay_registers_3_2_Im : _GEN_272; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_274 = 4'h3 == _GEN_270 ? input_delay_registers_3_3_Im : _GEN_273; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_275 = 4'h4 == _GEN_270 ? input_delay_registers_3_4_Im : _GEN_274; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_276 = 4'h5 == _GEN_270 ? input_delay_registers_3_5_Im : _GEN_275; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_277 = 4'h6 == _GEN_270 ? input_delay_registers_3_6_Im : _GEN_276; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_278 = 4'h7 == _GEN_270 ? input_delay_registers_3_7_Im : _GEN_277; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_279 = 4'h8 == _GEN_270 ? input_delay_registers_3_8_Im : _GEN_278; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_280 = 4'h9 == _GEN_270 ? input_delay_registers_3_9_Im : _GEN_279; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_281 = 4'ha == _GEN_270 ? input_delay_registers_3_10_Im : _GEN_280; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_282 = 4'hb == _GEN_270 ? input_delay_registers_3_11_Im : _GEN_281; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_284 = 4'h1 == _GEN_270 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_285 = 4'h2 == _GEN_270 ? input_delay_registers_3_2_Re : _GEN_284; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_286 = 4'h3 == _GEN_270 ? input_delay_registers_3_3_Re : _GEN_285; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_287 = 4'h4 == _GEN_270 ? input_delay_registers_3_4_Re : _GEN_286; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_288 = 4'h5 == _GEN_270 ? input_delay_registers_3_5_Re : _GEN_287; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_289 = 4'h6 == _GEN_270 ? input_delay_registers_3_6_Re : _GEN_288; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_290 = 4'h7 == _GEN_270 ? input_delay_registers_3_7_Re : _GEN_289; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_291 = 4'h8 == _GEN_270 ? input_delay_registers_3_8_Re : _GEN_290; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_292 = 4'h9 == _GEN_270 ? input_delay_registers_3_9_Re : _GEN_291; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_293 = 4'ha == _GEN_270 ? input_delay_registers_3_10_Re : _GEN_292; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_294 = 4'hb == _GEN_270 ? input_delay_registers_3_11_Re : _GEN_293; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_312 = 3'h1 == cnt ? 4'h7 : 4'h3; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_313 = 3'h2 == cnt ? 4'h3 : _GEN_312; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_314 = 3'h3 == cnt ? 4'h7 : _GEN_313; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_315 = 3'h4 == cnt ? 4'h3 : _GEN_314; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_316 = 3'h5 == cnt ? 4'h7 : _GEN_315; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_317 = 3'h6 == cnt ? 4'h3 : _GEN_316; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_318 = 3'h7 == cnt ? 4'h7 : _GEN_317; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_320 = 4'h1 == _GEN_318 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_321 = 4'h2 == _GEN_318 ? input_delay_registers_3_2_Im : _GEN_320; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_322 = 4'h3 == _GEN_318 ? input_delay_registers_3_3_Im : _GEN_321; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_323 = 4'h4 == _GEN_318 ? input_delay_registers_3_4_Im : _GEN_322; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_324 = 4'h5 == _GEN_318 ? input_delay_registers_3_5_Im : _GEN_323; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_325 = 4'h6 == _GEN_318 ? input_delay_registers_3_6_Im : _GEN_324; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_326 = 4'h7 == _GEN_318 ? input_delay_registers_3_7_Im : _GEN_325; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_327 = 4'h8 == _GEN_318 ? input_delay_registers_3_8_Im : _GEN_326; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_328 = 4'h9 == _GEN_318 ? input_delay_registers_3_9_Im : _GEN_327; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_329 = 4'ha == _GEN_318 ? input_delay_registers_3_10_Im : _GEN_328; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_330 = 4'hb == _GEN_318 ? input_delay_registers_3_11_Im : _GEN_329; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_332 = 4'h1 == _GEN_318 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_333 = 4'h2 == _GEN_318 ? input_delay_registers_3_2_Re : _GEN_332; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_334 = 4'h3 == _GEN_318 ? input_delay_registers_3_3_Re : _GEN_333; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_335 = 4'h4 == _GEN_318 ? input_delay_registers_3_4_Re : _GEN_334; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_336 = 4'h5 == _GEN_318 ? input_delay_registers_3_5_Re : _GEN_335; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_337 = 4'h6 == _GEN_318 ? input_delay_registers_3_6_Re : _GEN_336; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_338 = 4'h7 == _GEN_318 ? input_delay_registers_3_7_Re : _GEN_337; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_339 = 4'h8 == _GEN_318 ? input_delay_registers_3_8_Re : _GEN_338; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_340 = 4'h9 == _GEN_318 ? input_delay_registers_3_9_Re : _GEN_339; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_341 = 4'ha == _GEN_318 ? input_delay_registers_3_10_Re : _GEN_340; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_342 = 4'hb == _GEN_318 ? input_delay_registers_3_11_Re : _GEN_341; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_360 = 3'h1 == cnt ? 4'h0 : 4'hb; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_361 = 3'h2 == cnt ? 4'hb : _GEN_360; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_362 = 3'h3 == cnt ? 4'h0 : _GEN_361; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_363 = 3'h4 == cnt ? 4'hb : _GEN_362; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_364 = 3'h5 == cnt ? 4'h0 : _GEN_363; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_365 = 3'h6 == cnt ? 4'hb : _GEN_364; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_366 = 3'h7 == cnt ? 4'h0 : _GEN_365; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_368 = 4'h1 == _GEN_366 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_369 = 4'h2 == _GEN_366 ? input_delay_registers_3_2_Im : _GEN_368; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_370 = 4'h3 == _GEN_366 ? input_delay_registers_3_3_Im : _GEN_369; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_371 = 4'h4 == _GEN_366 ? input_delay_registers_3_4_Im : _GEN_370; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_372 = 4'h5 == _GEN_366 ? input_delay_registers_3_5_Im : _GEN_371; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_373 = 4'h6 == _GEN_366 ? input_delay_registers_3_6_Im : _GEN_372; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_374 = 4'h7 == _GEN_366 ? input_delay_registers_3_7_Im : _GEN_373; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_375 = 4'h8 == _GEN_366 ? input_delay_registers_3_8_Im : _GEN_374; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_376 = 4'h9 == _GEN_366 ? input_delay_registers_3_9_Im : _GEN_375; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_377 = 4'ha == _GEN_366 ? input_delay_registers_3_10_Im : _GEN_376; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_378 = 4'hb == _GEN_366 ? input_delay_registers_3_11_Im : _GEN_377; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_380 = 4'h1 == _GEN_366 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_381 = 4'h2 == _GEN_366 ? input_delay_registers_3_2_Re : _GEN_380; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_382 = 4'h3 == _GEN_366 ? input_delay_registers_3_3_Re : _GEN_381; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_383 = 4'h4 == _GEN_366 ? input_delay_registers_3_4_Re : _GEN_382; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_384 = 4'h5 == _GEN_366 ? input_delay_registers_3_5_Re : _GEN_383; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_385 = 4'h6 == _GEN_366 ? input_delay_registers_3_6_Re : _GEN_384; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_386 = 4'h7 == _GEN_366 ? input_delay_registers_3_7_Re : _GEN_385; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_387 = 4'h8 == _GEN_366 ? input_delay_registers_3_8_Re : _GEN_386; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_388 = 4'h9 == _GEN_366 ? input_delay_registers_3_9_Re : _GEN_387; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_389 = 4'ha == _GEN_366 ? input_delay_registers_3_10_Re : _GEN_388; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_390 = 4'hb == _GEN_366 ? input_delay_registers_3_11_Re : _GEN_389; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_400 = 3'h1 == cnt ? 4'h1 : 4'h0; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_401 = 3'h2 == cnt ? 4'h3 : _GEN_400; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_402 = 3'h3 == cnt ? 4'h4 : _GEN_401; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_403 = 3'h4 == cnt ? 4'h6 : _GEN_402; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_404 = 3'h5 == cnt ? 4'h7 : _GEN_403; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_405 = 3'h6 == cnt ? 4'h9 : _GEN_404; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_406 = 3'h7 == cnt ? 4'ha : _GEN_405; // @[FFTDesigns.scala 2978:{55,55}]
  wire [4:0] _GEN_1052 = {{1'd0}, _GEN_406}; // @[FFTDesigns.scala 2978:55]
  wire [4:0] _M0_4_in_waddr_0_T_2 = _GEN_1052 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2978:55]
  wire [3:0] _GEN_408 = 3'h1 == cnt ? 4'h0 : 4'h4; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_409 = 3'h2 == cnt ? 4'h4 : _GEN_408; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_410 = 3'h3 == cnt ? 4'h0 : _GEN_409; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_411 = 3'h4 == cnt ? 4'h4 : _GEN_410; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_412 = 3'h5 == cnt ? 4'h0 : _GEN_411; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_413 = 3'h6 == cnt ? 4'h4 : _GEN_412; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_414 = 3'h7 == cnt ? 4'h0 : _GEN_413; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_416 = 4'h1 == _GEN_414 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_417 = 4'h2 == _GEN_414 ? input_delay_registers_3_2_Im : _GEN_416; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_418 = 4'h3 == _GEN_414 ? input_delay_registers_3_3_Im : _GEN_417; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_419 = 4'h4 == _GEN_414 ? input_delay_registers_3_4_Im : _GEN_418; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_420 = 4'h5 == _GEN_414 ? input_delay_registers_3_5_Im : _GEN_419; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_421 = 4'h6 == _GEN_414 ? input_delay_registers_3_6_Im : _GEN_420; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_422 = 4'h7 == _GEN_414 ? input_delay_registers_3_7_Im : _GEN_421; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_423 = 4'h8 == _GEN_414 ? input_delay_registers_3_8_Im : _GEN_422; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_424 = 4'h9 == _GEN_414 ? input_delay_registers_3_9_Im : _GEN_423; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_425 = 4'ha == _GEN_414 ? input_delay_registers_3_10_Im : _GEN_424; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_426 = 4'hb == _GEN_414 ? input_delay_registers_3_11_Im : _GEN_425; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_428 = 4'h1 == _GEN_414 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_429 = 4'h2 == _GEN_414 ? input_delay_registers_3_2_Re : _GEN_428; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_430 = 4'h3 == _GEN_414 ? input_delay_registers_3_3_Re : _GEN_429; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_431 = 4'h4 == _GEN_414 ? input_delay_registers_3_4_Re : _GEN_430; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_432 = 4'h5 == _GEN_414 ? input_delay_registers_3_5_Re : _GEN_431; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_433 = 4'h6 == _GEN_414 ? input_delay_registers_3_6_Re : _GEN_432; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_434 = 4'h7 == _GEN_414 ? input_delay_registers_3_7_Re : _GEN_433; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_435 = 4'h8 == _GEN_414 ? input_delay_registers_3_8_Re : _GEN_434; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_436 = 4'h9 == _GEN_414 ? input_delay_registers_3_9_Re : _GEN_435; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_437 = 4'ha == _GEN_414 ? input_delay_registers_3_10_Re : _GEN_436; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_438 = 4'hb == _GEN_414 ? input_delay_registers_3_11_Re : _GEN_437; // @[FFTDesigns.scala 2979:{32,32}]
  wire  _GEN_441 = 3'h2 == cnt ? 1'h0 : 3'h1 == cnt; // @[FFTDesigns.scala 2977:{27,27}]
  wire  _GEN_443 = 3'h4 == cnt ? 1'h0 : 3'h3 == cnt | _GEN_441; // @[FFTDesigns.scala 2977:{27,27}]
  wire  _GEN_445 = 3'h6 == cnt ? 1'h0 : 3'h5 == cnt | _GEN_443; // @[FFTDesigns.scala 2977:{27,27}]
  wire [3:0] _GEN_449 = 3'h2 == cnt ? 4'h0 : _GEN_16; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_450 = 3'h3 == cnt ? 4'h5 : _GEN_449; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_451 = 3'h4 == cnt ? 4'h0 : _GEN_450; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_452 = 3'h5 == cnt ? 4'h8 : _GEN_451; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_453 = 3'h6 == cnt ? 4'h0 : _GEN_452; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_454 = 3'h7 == cnt ? 4'hb : _GEN_453; // @[FFTDesigns.scala 2978:{55,55}]
  wire [4:0] _GEN_1056 = {{1'd0}, _GEN_454}; // @[FFTDesigns.scala 2978:55]
  wire [4:0] _M0_4_in_waddr_1_T_2 = _GEN_1056 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2978:55]
  wire [3:0] _GEN_456 = 3'h1 == cnt ? 4'h8 : 4'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_457 = 3'h2 == cnt ? 4'h0 : _GEN_456; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_458 = 3'h3 == cnt ? 4'h8 : _GEN_457; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_459 = 3'h4 == cnt ? 4'h0 : _GEN_458; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_460 = 3'h5 == cnt ? 4'h8 : _GEN_459; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_461 = 3'h6 == cnt ? 4'h0 : _GEN_460; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_462 = 3'h7 == cnt ? 4'h8 : _GEN_461; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_464 = 4'h1 == _GEN_462 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_465 = 4'h2 == _GEN_462 ? input_delay_registers_3_2_Im : _GEN_464; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_466 = 4'h3 == _GEN_462 ? input_delay_registers_3_3_Im : _GEN_465; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_467 = 4'h4 == _GEN_462 ? input_delay_registers_3_4_Im : _GEN_466; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_468 = 4'h5 == _GEN_462 ? input_delay_registers_3_5_Im : _GEN_467; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_469 = 4'h6 == _GEN_462 ? input_delay_registers_3_6_Im : _GEN_468; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_470 = 4'h7 == _GEN_462 ? input_delay_registers_3_7_Im : _GEN_469; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_471 = 4'h8 == _GEN_462 ? input_delay_registers_3_8_Im : _GEN_470; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_472 = 4'h9 == _GEN_462 ? input_delay_registers_3_9_Im : _GEN_471; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_473 = 4'ha == _GEN_462 ? input_delay_registers_3_10_Im : _GEN_472; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_474 = 4'hb == _GEN_462 ? input_delay_registers_3_11_Im : _GEN_473; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_476 = 4'h1 == _GEN_462 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_477 = 4'h2 == _GEN_462 ? input_delay_registers_3_2_Re : _GEN_476; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_478 = 4'h3 == _GEN_462 ? input_delay_registers_3_3_Re : _GEN_477; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_479 = 4'h4 == _GEN_462 ? input_delay_registers_3_4_Re : _GEN_478; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_480 = 4'h5 == _GEN_462 ? input_delay_registers_3_5_Re : _GEN_479; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_481 = 4'h6 == _GEN_462 ? input_delay_registers_3_6_Re : _GEN_480; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_482 = 4'h7 == _GEN_462 ? input_delay_registers_3_7_Re : _GEN_481; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_483 = 4'h8 == _GEN_462 ? input_delay_registers_3_8_Re : _GEN_482; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_484 = 4'h9 == _GEN_462 ? input_delay_registers_3_9_Re : _GEN_483; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_485 = 4'ha == _GEN_462 ? input_delay_registers_3_10_Re : _GEN_484; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_486 = 4'hb == _GEN_462 ? input_delay_registers_3_11_Re : _GEN_485; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_504 = 3'h1 == cnt ? 4'h1 : 4'h5; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_505 = 3'h2 == cnt ? 4'h5 : _GEN_504; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_506 = 3'h3 == cnt ? 4'h1 : _GEN_505; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_507 = 3'h4 == cnt ? 4'h5 : _GEN_506; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_508 = 3'h5 == cnt ? 4'h1 : _GEN_507; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_509 = 3'h6 == cnt ? 4'h5 : _GEN_508; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_510 = 3'h7 == cnt ? 4'h1 : _GEN_509; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_512 = 4'h1 == _GEN_510 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_513 = 4'h2 == _GEN_510 ? input_delay_registers_3_2_Im : _GEN_512; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_514 = 4'h3 == _GEN_510 ? input_delay_registers_3_3_Im : _GEN_513; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_515 = 4'h4 == _GEN_510 ? input_delay_registers_3_4_Im : _GEN_514; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_516 = 4'h5 == _GEN_510 ? input_delay_registers_3_5_Im : _GEN_515; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_517 = 4'h6 == _GEN_510 ? input_delay_registers_3_6_Im : _GEN_516; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_518 = 4'h7 == _GEN_510 ? input_delay_registers_3_7_Im : _GEN_517; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_519 = 4'h8 == _GEN_510 ? input_delay_registers_3_8_Im : _GEN_518; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_520 = 4'h9 == _GEN_510 ? input_delay_registers_3_9_Im : _GEN_519; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_521 = 4'ha == _GEN_510 ? input_delay_registers_3_10_Im : _GEN_520; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_522 = 4'hb == _GEN_510 ? input_delay_registers_3_11_Im : _GEN_521; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_524 = 4'h1 == _GEN_510 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_525 = 4'h2 == _GEN_510 ? input_delay_registers_3_2_Re : _GEN_524; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_526 = 4'h3 == _GEN_510 ? input_delay_registers_3_3_Re : _GEN_525; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_527 = 4'h4 == _GEN_510 ? input_delay_registers_3_4_Re : _GEN_526; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_528 = 4'h5 == _GEN_510 ? input_delay_registers_3_5_Re : _GEN_527; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_529 = 4'h6 == _GEN_510 ? input_delay_registers_3_6_Re : _GEN_528; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_530 = 4'h7 == _GEN_510 ? input_delay_registers_3_7_Re : _GEN_529; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_531 = 4'h8 == _GEN_510 ? input_delay_registers_3_8_Re : _GEN_530; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_532 = 4'h9 == _GEN_510 ? input_delay_registers_3_9_Re : _GEN_531; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_533 = 4'ha == _GEN_510 ? input_delay_registers_3_10_Re : _GEN_532; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_534 = 4'hb == _GEN_510 ? input_delay_registers_3_11_Re : _GEN_533; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_552 = 3'h1 == cnt ? 4'h9 : 4'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_553 = 3'h2 == cnt ? 4'h0 : _GEN_552; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_554 = 3'h3 == cnt ? 4'h9 : _GEN_553; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_555 = 3'h4 == cnt ? 4'h0 : _GEN_554; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_556 = 3'h5 == cnt ? 4'h9 : _GEN_555; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_557 = 3'h6 == cnt ? 4'h0 : _GEN_556; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_558 = 3'h7 == cnt ? 4'h9 : _GEN_557; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_560 = 4'h1 == _GEN_558 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_561 = 4'h2 == _GEN_558 ? input_delay_registers_3_2_Im : _GEN_560; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_562 = 4'h3 == _GEN_558 ? input_delay_registers_3_3_Im : _GEN_561; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_563 = 4'h4 == _GEN_558 ? input_delay_registers_3_4_Im : _GEN_562; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_564 = 4'h5 == _GEN_558 ? input_delay_registers_3_5_Im : _GEN_563; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_565 = 4'h6 == _GEN_558 ? input_delay_registers_3_6_Im : _GEN_564; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_566 = 4'h7 == _GEN_558 ? input_delay_registers_3_7_Im : _GEN_565; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_567 = 4'h8 == _GEN_558 ? input_delay_registers_3_8_Im : _GEN_566; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_568 = 4'h9 == _GEN_558 ? input_delay_registers_3_9_Im : _GEN_567; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_569 = 4'ha == _GEN_558 ? input_delay_registers_3_10_Im : _GEN_568; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_570 = 4'hb == _GEN_558 ? input_delay_registers_3_11_Im : _GEN_569; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_572 = 4'h1 == _GEN_558 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_573 = 4'h2 == _GEN_558 ? input_delay_registers_3_2_Re : _GEN_572; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_574 = 4'h3 == _GEN_558 ? input_delay_registers_3_3_Re : _GEN_573; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_575 = 4'h4 == _GEN_558 ? input_delay_registers_3_4_Re : _GEN_574; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_576 = 4'h5 == _GEN_558 ? input_delay_registers_3_5_Re : _GEN_575; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_577 = 4'h6 == _GEN_558 ? input_delay_registers_3_6_Re : _GEN_576; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_578 = 4'h7 == _GEN_558 ? input_delay_registers_3_7_Re : _GEN_577; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_579 = 4'h8 == _GEN_558 ? input_delay_registers_3_8_Re : _GEN_578; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_580 = 4'h9 == _GEN_558 ? input_delay_registers_3_9_Re : _GEN_579; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_581 = 4'ha == _GEN_558 ? input_delay_registers_3_10_Re : _GEN_580; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_582 = 4'hb == _GEN_558 ? input_delay_registers_3_11_Re : _GEN_581; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_600 = 3'h1 == cnt ? 4'h2 : 4'h6; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_601 = 3'h2 == cnt ? 4'h6 : _GEN_600; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_602 = 3'h3 == cnt ? 4'h2 : _GEN_601; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_603 = 3'h4 == cnt ? 4'h6 : _GEN_602; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_604 = 3'h5 == cnt ? 4'h2 : _GEN_603; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_605 = 3'h6 == cnt ? 4'h6 : _GEN_604; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_606 = 3'h7 == cnt ? 4'h2 : _GEN_605; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_608 = 4'h1 == _GEN_606 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_609 = 4'h2 == _GEN_606 ? input_delay_registers_3_2_Im : _GEN_608; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_610 = 4'h3 == _GEN_606 ? input_delay_registers_3_3_Im : _GEN_609; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_611 = 4'h4 == _GEN_606 ? input_delay_registers_3_4_Im : _GEN_610; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_612 = 4'h5 == _GEN_606 ? input_delay_registers_3_5_Im : _GEN_611; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_613 = 4'h6 == _GEN_606 ? input_delay_registers_3_6_Im : _GEN_612; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_614 = 4'h7 == _GEN_606 ? input_delay_registers_3_7_Im : _GEN_613; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_615 = 4'h8 == _GEN_606 ? input_delay_registers_3_8_Im : _GEN_614; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_616 = 4'h9 == _GEN_606 ? input_delay_registers_3_9_Im : _GEN_615; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_617 = 4'ha == _GEN_606 ? input_delay_registers_3_10_Im : _GEN_616; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_618 = 4'hb == _GEN_606 ? input_delay_registers_3_11_Im : _GEN_617; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_620 = 4'h1 == _GEN_606 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_621 = 4'h2 == _GEN_606 ? input_delay_registers_3_2_Re : _GEN_620; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_622 = 4'h3 == _GEN_606 ? input_delay_registers_3_3_Re : _GEN_621; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_623 = 4'h4 == _GEN_606 ? input_delay_registers_3_4_Re : _GEN_622; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_624 = 4'h5 == _GEN_606 ? input_delay_registers_3_5_Re : _GEN_623; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_625 = 4'h6 == _GEN_606 ? input_delay_registers_3_6_Re : _GEN_624; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_626 = 4'h7 == _GEN_606 ? input_delay_registers_3_7_Re : _GEN_625; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_627 = 4'h8 == _GEN_606 ? input_delay_registers_3_8_Re : _GEN_626; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_628 = 4'h9 == _GEN_606 ? input_delay_registers_3_9_Re : _GEN_627; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_629 = 4'ha == _GEN_606 ? input_delay_registers_3_10_Re : _GEN_628; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_630 = 4'hb == _GEN_606 ? input_delay_registers_3_11_Re : _GEN_629; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_648 = 3'h1 == cnt ? 4'ha : 4'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_649 = 3'h2 == cnt ? 4'h0 : _GEN_648; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_650 = 3'h3 == cnt ? 4'ha : _GEN_649; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_651 = 3'h4 == cnt ? 4'h0 : _GEN_650; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_652 = 3'h5 == cnt ? 4'ha : _GEN_651; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_653 = 3'h6 == cnt ? 4'h0 : _GEN_652; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_654 = 3'h7 == cnt ? 4'ha : _GEN_653; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_656 = 4'h1 == _GEN_654 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_657 = 4'h2 == _GEN_654 ? input_delay_registers_3_2_Im : _GEN_656; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_658 = 4'h3 == _GEN_654 ? input_delay_registers_3_3_Im : _GEN_657; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_659 = 4'h4 == _GEN_654 ? input_delay_registers_3_4_Im : _GEN_658; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_660 = 4'h5 == _GEN_654 ? input_delay_registers_3_5_Im : _GEN_659; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_661 = 4'h6 == _GEN_654 ? input_delay_registers_3_6_Im : _GEN_660; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_662 = 4'h7 == _GEN_654 ? input_delay_registers_3_7_Im : _GEN_661; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_663 = 4'h8 == _GEN_654 ? input_delay_registers_3_8_Im : _GEN_662; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_664 = 4'h9 == _GEN_654 ? input_delay_registers_3_9_Im : _GEN_663; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_665 = 4'ha == _GEN_654 ? input_delay_registers_3_10_Im : _GEN_664; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_666 = 4'hb == _GEN_654 ? input_delay_registers_3_11_Im : _GEN_665; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_668 = 4'h1 == _GEN_654 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_669 = 4'h2 == _GEN_654 ? input_delay_registers_3_2_Re : _GEN_668; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_670 = 4'h3 == _GEN_654 ? input_delay_registers_3_3_Re : _GEN_669; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_671 = 4'h4 == _GEN_654 ? input_delay_registers_3_4_Re : _GEN_670; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_672 = 4'h5 == _GEN_654 ? input_delay_registers_3_5_Re : _GEN_671; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_673 = 4'h6 == _GEN_654 ? input_delay_registers_3_6_Re : _GEN_672; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_674 = 4'h7 == _GEN_654 ? input_delay_registers_3_7_Re : _GEN_673; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_675 = 4'h8 == _GEN_654 ? input_delay_registers_3_8_Re : _GEN_674; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_676 = 4'h9 == _GEN_654 ? input_delay_registers_3_9_Re : _GEN_675; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_677 = 4'ha == _GEN_654 ? input_delay_registers_3_10_Re : _GEN_676; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_678 = 4'hb == _GEN_654 ? input_delay_registers_3_11_Re : _GEN_677; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_696 = 3'h1 == cnt ? 4'h3 : 4'h7; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_697 = 3'h2 == cnt ? 4'h7 : _GEN_696; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_698 = 3'h3 == cnt ? 4'h3 : _GEN_697; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_699 = 3'h4 == cnt ? 4'h7 : _GEN_698; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_700 = 3'h5 == cnt ? 4'h3 : _GEN_699; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_701 = 3'h6 == cnt ? 4'h7 : _GEN_700; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_702 = 3'h7 == cnt ? 4'h3 : _GEN_701; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_704 = 4'h1 == _GEN_702 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_705 = 4'h2 == _GEN_702 ? input_delay_registers_3_2_Im : _GEN_704; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_706 = 4'h3 == _GEN_702 ? input_delay_registers_3_3_Im : _GEN_705; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_707 = 4'h4 == _GEN_702 ? input_delay_registers_3_4_Im : _GEN_706; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_708 = 4'h5 == _GEN_702 ? input_delay_registers_3_5_Im : _GEN_707; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_709 = 4'h6 == _GEN_702 ? input_delay_registers_3_6_Im : _GEN_708; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_710 = 4'h7 == _GEN_702 ? input_delay_registers_3_7_Im : _GEN_709; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_711 = 4'h8 == _GEN_702 ? input_delay_registers_3_8_Im : _GEN_710; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_712 = 4'h9 == _GEN_702 ? input_delay_registers_3_9_Im : _GEN_711; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_713 = 4'ha == _GEN_702 ? input_delay_registers_3_10_Im : _GEN_712; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_714 = 4'hb == _GEN_702 ? input_delay_registers_3_11_Im : _GEN_713; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_716 = 4'h1 == _GEN_702 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_717 = 4'h2 == _GEN_702 ? input_delay_registers_3_2_Re : _GEN_716; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_718 = 4'h3 == _GEN_702 ? input_delay_registers_3_3_Re : _GEN_717; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_719 = 4'h4 == _GEN_702 ? input_delay_registers_3_4_Re : _GEN_718; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_720 = 4'h5 == _GEN_702 ? input_delay_registers_3_5_Re : _GEN_719; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_721 = 4'h6 == _GEN_702 ? input_delay_registers_3_6_Re : _GEN_720; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_722 = 4'h7 == _GEN_702 ? input_delay_registers_3_7_Re : _GEN_721; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_723 = 4'h8 == _GEN_702 ? input_delay_registers_3_8_Re : _GEN_722; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_724 = 4'h9 == _GEN_702 ? input_delay_registers_3_9_Re : _GEN_723; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_725 = 4'ha == _GEN_702 ? input_delay_registers_3_10_Re : _GEN_724; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_726 = 4'hb == _GEN_702 ? input_delay_registers_3_11_Re : _GEN_725; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_744 = 3'h1 == cnt ? 4'hb : 4'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_745 = 3'h2 == cnt ? 4'h0 : _GEN_744; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_746 = 3'h3 == cnt ? 4'hb : _GEN_745; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_747 = 3'h4 == cnt ? 4'h0 : _GEN_746; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_748 = 3'h5 == cnt ? 4'hb : _GEN_747; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_749 = 3'h6 == cnt ? 4'h0 : _GEN_748; // @[FFTDesigns.scala 2979:{32,32}]
  wire [3:0] _GEN_750 = 3'h7 == cnt ? 4'hb : _GEN_749; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_752 = 4'h1 == _GEN_750 ? input_delay_registers_3_1_Im : input_delay_registers_3_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_753 = 4'h2 == _GEN_750 ? input_delay_registers_3_2_Im : _GEN_752; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_754 = 4'h3 == _GEN_750 ? input_delay_registers_3_3_Im : _GEN_753; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_755 = 4'h4 == _GEN_750 ? input_delay_registers_3_4_Im : _GEN_754; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_756 = 4'h5 == _GEN_750 ? input_delay_registers_3_5_Im : _GEN_755; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_757 = 4'h6 == _GEN_750 ? input_delay_registers_3_6_Im : _GEN_756; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_758 = 4'h7 == _GEN_750 ? input_delay_registers_3_7_Im : _GEN_757; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_759 = 4'h8 == _GEN_750 ? input_delay_registers_3_8_Im : _GEN_758; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_760 = 4'h9 == _GEN_750 ? input_delay_registers_3_9_Im : _GEN_759; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_761 = 4'ha == _GEN_750 ? input_delay_registers_3_10_Im : _GEN_760; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_762 = 4'hb == _GEN_750 ? input_delay_registers_3_11_Im : _GEN_761; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_764 = 4'h1 == _GEN_750 ? input_delay_registers_3_1_Re : input_delay_registers_3_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_765 = 4'h2 == _GEN_750 ? input_delay_registers_3_2_Re : _GEN_764; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_766 = 4'h3 == _GEN_750 ? input_delay_registers_3_3_Re : _GEN_765; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_767 = 4'h4 == _GEN_750 ? input_delay_registers_3_4_Re : _GEN_766; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_768 = 4'h5 == _GEN_750 ? input_delay_registers_3_5_Re : _GEN_767; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_769 = 4'h6 == _GEN_750 ? input_delay_registers_3_6_Re : _GEN_768; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_770 = 4'h7 == _GEN_750 ? input_delay_registers_3_7_Re : _GEN_769; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_771 = 4'h8 == _GEN_750 ? input_delay_registers_3_8_Re : _GEN_770; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_772 = 4'h9 == _GEN_750 ? input_delay_registers_3_9_Re : _GEN_771; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_773 = 4'ha == _GEN_750 ? input_delay_registers_3_10_Re : _GEN_772; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_774 = 4'hb == _GEN_750 ? input_delay_registers_3_11_Re : _GEN_773; // @[FFTDesigns.scala 2979:{32,32}]
  RAM_Block_mw RAM_Block_mw ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_clock),
    .io_in_raddr(RAM_Block_mw_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_io_in_data_1_Im),
    .io_re(RAM_Block_mw_io_re),
    .io_wr_0(RAM_Block_mw_io_wr_0),
    .io_wr_1(RAM_Block_mw_io_wr_1),
    .io_en(RAM_Block_mw_io_en),
    .io_out_data_Re(RAM_Block_mw_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_1 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_1_clock),
    .io_in_raddr(RAM_Block_mw_1_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_1_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_1_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_1_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_1_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_1_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_1_io_in_data_1_Im),
    .io_re(RAM_Block_mw_1_io_re),
    .io_wr_0(RAM_Block_mw_1_io_wr_0),
    .io_wr_1(RAM_Block_mw_1_io_wr_1),
    .io_en(RAM_Block_mw_1_io_en),
    .io_out_data_Re(RAM_Block_mw_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_1_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_2 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_2_clock),
    .io_in_raddr(RAM_Block_mw_2_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_2_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_2_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_2_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_2_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_2_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_2_io_in_data_1_Im),
    .io_re(RAM_Block_mw_2_io_re),
    .io_wr_0(RAM_Block_mw_2_io_wr_0),
    .io_wr_1(RAM_Block_mw_2_io_wr_1),
    .io_en(RAM_Block_mw_2_io_en),
    .io_out_data_Re(RAM_Block_mw_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_2_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_3 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_3_clock),
    .io_in_raddr(RAM_Block_mw_3_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_3_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_3_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_3_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_3_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_3_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_3_io_in_data_1_Im),
    .io_re(RAM_Block_mw_3_io_re),
    .io_wr_0(RAM_Block_mw_3_io_wr_0),
    .io_wr_1(RAM_Block_mw_3_io_wr_1),
    .io_en(RAM_Block_mw_3_io_en),
    .io_out_data_Re(RAM_Block_mw_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_3_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_4 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_4_clock),
    .io_in_raddr(RAM_Block_mw_4_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_4_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_4_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_4_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_4_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_4_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_4_io_in_data_1_Im),
    .io_re(RAM_Block_mw_4_io_re),
    .io_wr_0(RAM_Block_mw_4_io_wr_0),
    .io_wr_1(RAM_Block_mw_4_io_wr_1),
    .io_en(RAM_Block_mw_4_io_en),
    .io_out_data_Re(RAM_Block_mw_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_4_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_5 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_5_clock),
    .io_in_raddr(RAM_Block_mw_5_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_5_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_5_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_5_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_5_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_5_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_5_io_in_data_1_Im),
    .io_re(RAM_Block_mw_5_io_re),
    .io_wr_0(RAM_Block_mw_5_io_wr_0),
    .io_wr_1(RAM_Block_mw_5_io_wr_1),
    .io_en(RAM_Block_mw_5_io_en),
    .io_out_data_Re(RAM_Block_mw_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_5_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_6 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_6_clock),
    .io_in_raddr(RAM_Block_mw_6_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_6_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_6_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_6_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_6_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_6_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_6_io_in_data_1_Im),
    .io_re(RAM_Block_mw_6_io_re),
    .io_wr_0(RAM_Block_mw_6_io_wr_0),
    .io_wr_1(RAM_Block_mw_6_io_wr_1),
    .io_en(RAM_Block_mw_6_io_en),
    .io_out_data_Re(RAM_Block_mw_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_6_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_7 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_7_clock),
    .io_in_raddr(RAM_Block_mw_7_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_7_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_7_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_7_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_7_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_7_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_7_io_in_data_1_Im),
    .io_re(RAM_Block_mw_7_io_re),
    .io_wr_0(RAM_Block_mw_7_io_wr_0),
    .io_wr_1(RAM_Block_mw_7_io_wr_1),
    .io_en(RAM_Block_mw_7_io_en),
    .io_out_data_Re(RAM_Block_mw_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_7_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_1 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_2 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_3 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_4 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_5 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_6 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block_96 RAM_Block_7 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  PermutationModuleStreamed PermutationModuleStreamed ( // @[FFTDesigns.scala 2907:28]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im)
  );
  M0_Config_ROM_6 M0_Config_ROM ( // @[FFTDesigns.scala 2908:29]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7)
  );
  M1_Config_ROM_6 M1_Config_ROM ( // @[FFTDesigns.scala 2909:29]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7)
  );
  Streaming_Permute_Config_6 Streaming_Permute_Config ( // @[FFTDesigns.scala 2910:31]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6)
  );
  assign io_out_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign RAM_Block_mw_clock = clock;
  assign RAM_Block_mw_io_in_raddr = M0_0_re ? _M0_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_io_in_data_0_Re = M0_0_re ? _GEN_54 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_io_in_data_0_Im = M0_0_re ? _GEN_42 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_io_in_data_1_Re = M0_0_re ? _GEN_102 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_io_in_data_1_Im = M0_0_re ? _GEN_90 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_io_wr_1 = M0_0_re & _GEN_62; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_1_clock = clock;
  assign RAM_Block_mw_1_io_in_raddr = M0_0_re ? _M0_1_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_1_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_1_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_1_io_in_data_0_Re = M0_0_re ? _GEN_150 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_1_io_in_data_0_Im = M0_0_re ? _GEN_138 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_1_io_in_data_1_Re = M0_0_re ? _GEN_198 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_1_io_in_data_1_Im = M0_0_re ? _GEN_186 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_1_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_1_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_1_io_wr_1 = M0_0_re & _GEN_62; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_1_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_2_clock = clock;
  assign RAM_Block_mw_2_io_in_raddr = M0_0_re ? _M0_2_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_2_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_2_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_2_io_in_data_0_Re = M0_0_re ? _GEN_246 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_2_io_in_data_0_Im = M0_0_re ? _GEN_234 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_2_io_in_data_1_Re = M0_0_re ? _GEN_294 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_2_io_in_data_1_Im = M0_0_re ? _GEN_282 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_2_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_2_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_2_io_wr_1 = M0_0_re & _GEN_62; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_2_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_3_clock = clock;
  assign RAM_Block_mw_3_io_in_raddr = M0_0_re ? _M0_3_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_3_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_3_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_3_io_in_data_0_Re = M0_0_re ? _GEN_342 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_3_io_in_data_0_Im = M0_0_re ? _GEN_330 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_3_io_in_data_1_Re = M0_0_re ? _GEN_390 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_3_io_in_data_1_Im = M0_0_re ? _GEN_378 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_3_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_3_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_3_io_wr_1 = M0_0_re & _GEN_62; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_3_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_4_clock = clock;
  assign RAM_Block_mw_4_io_in_raddr = M0_0_re ? _M0_4_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_4_io_in_waddr_0 = M0_0_re ? _M0_4_in_waddr_0_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_4_io_in_waddr_1 = M0_0_re ? _M0_4_in_waddr_1_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_4_io_in_data_0_Re = M0_0_re ? _GEN_438 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_4_io_in_data_0_Im = M0_0_re ? _GEN_426 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_4_io_in_data_1_Re = M0_0_re ? _GEN_486 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_4_io_in_data_1_Im = M0_0_re ? _GEN_474 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_4_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_4_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_4_io_wr_1 = M0_0_re & (3'h7 == cnt | _GEN_445); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_4_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_5_clock = clock;
  assign RAM_Block_mw_5_io_in_raddr = M0_0_re ? _M0_5_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_5_io_in_waddr_0 = M0_0_re ? _M0_4_in_waddr_0_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_5_io_in_waddr_1 = M0_0_re ? _M0_4_in_waddr_1_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_5_io_in_data_0_Re = M0_0_re ? _GEN_534 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_5_io_in_data_0_Im = M0_0_re ? _GEN_522 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_5_io_in_data_1_Re = M0_0_re ? _GEN_582 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_5_io_in_data_1_Im = M0_0_re ? _GEN_570 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_5_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_5_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_5_io_wr_1 = M0_0_re & (3'h7 == cnt | _GEN_445); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_5_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_6_clock = clock;
  assign RAM_Block_mw_6_io_in_raddr = M0_0_re ? _M0_6_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_6_io_in_waddr_0 = M0_0_re ? _M0_4_in_waddr_0_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_6_io_in_waddr_1 = M0_0_re ? _M0_4_in_waddr_1_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_6_io_in_data_0_Re = M0_0_re ? _GEN_630 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_6_io_in_data_0_Im = M0_0_re ? _GEN_618 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_6_io_in_data_1_Re = M0_0_re ? _GEN_678 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_6_io_in_data_1_Im = M0_0_re ? _GEN_666 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_6_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_6_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_6_io_wr_1 = M0_0_re & (3'h7 == cnt | _GEN_445); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_6_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_7_clock = clock;
  assign RAM_Block_mw_7_io_in_raddr = M0_0_re ? _M0_7_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_7_io_in_waddr_0 = M0_0_re ? _M0_4_in_waddr_0_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_7_io_in_waddr_1 = M0_0_re ? _M0_4_in_waddr_1_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_7_io_in_data_0_Re = M0_0_re ? _GEN_726 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_7_io_in_data_0_Im = M0_0_re ? _GEN_714 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_7_io_in_data_1_Re = M0_0_re ? _GEN_774 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_7_io_in_data_1_Im = M0_0_re ? _GEN_762 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_7_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_7_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_7_io_wr_1 = M0_0_re & (3'h7 == cnt | _GEN_445); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_7_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_io_in_waddr = M0_0_re ? _M1_0_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_1_io_in_waddr = M0_0_re ? _M1_1_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_1_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_1_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_1_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_2_io_in_waddr = M0_0_re ? _M1_2_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_2_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_2_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_2_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_3_io_in_waddr = M0_0_re ? _M1_3_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_3_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_3_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_3_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_4_io_in_waddr = M0_0_re ? _M1_4_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_4_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_4_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_4_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_5_io_in_waddr = M0_0_re ? _M1_5_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_5_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_5_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_5_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_6_io_in_waddr = M0_0_re ? _M1_6_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_6_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_6_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_6_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 5'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_7_io_in_waddr = M0_0_re ? _M1_7_in_waddr_T_2 : 5'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_7_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_7_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_7_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_mw_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_mw_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_mw_1_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_mw_1_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_mw_2_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_mw_2_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_mw_3_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_mw_3_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_mw_4_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_mw_4_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_mw_5_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_mw_5_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_mw_6_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_mw_6_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_mw_7_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_mw_7_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign M0_Config_ROM_io_in_cnt = cnt2; // @[FFTDesigns.scala 3021:24]
  assign M1_Config_ROM_io_in_cnt = cnt2; // @[FFTDesigns.scala 3022:24]
  assign Streaming_Permute_Config_io_in_cnt = cnt2; // @[FFTDesigns.scala 3023:26]
  always @(posedge clock) begin
    offset_switch <= M0_0_re & _GEN_6; // @[FFTDesigns.scala 2914:33 3017:23]
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_0_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_0_Re <= io_in_0_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_0_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_0_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_0_Im <= io_in_0_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_0_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_1_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_1_Re <= io_in_1_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_1_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_1_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_1_Im <= io_in_1_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_1_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_2_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_2_Re <= io_in_2_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_2_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_2_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_2_Im <= io_in_2_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_2_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_3_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_3_Re <= io_in_3_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_3_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_3_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_3_Im <= io_in_3_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_3_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_4_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_4_Re <= io_in_4_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_4_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_4_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_4_Im <= io_in_4_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_4_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_5_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_5_Re <= io_in_5_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_5_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_5_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_5_Im <= io_in_5_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_5_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_6_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_6_Re <= io_in_6_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_6_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_6_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_6_Im <= io_in_6_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_6_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_7_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_7_Re <= io_in_7_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_7_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_7_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_7_Im <= io_in_7_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_7_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_8_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_8_Re <= io_in_8_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_8_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_8_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_8_Im <= io_in_8_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_8_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_9_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_9_Re <= io_in_9_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_9_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_9_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_9_Im <= io_in_9_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_9_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_10_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_10_Re <= io_in_10_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_10_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_10_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_10_Im <= io_in_10_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_10_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_11_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_11_Re <= io_in_11_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_11_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_11_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_11_Im <= io_in_11_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_11_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_0_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_0_Re <= input_delay_registers_0_0_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_0_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_0_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_0_Im <= input_delay_registers_0_0_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_0_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_1_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_1_Re <= input_delay_registers_0_1_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_1_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_1_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_1_Im <= input_delay_registers_0_1_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_1_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_2_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_2_Re <= input_delay_registers_0_2_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_2_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_2_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_2_Im <= input_delay_registers_0_2_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_2_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_3_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_3_Re <= input_delay_registers_0_3_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_3_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_3_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_3_Im <= input_delay_registers_0_3_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_3_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_4_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_4_Re <= input_delay_registers_0_4_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_4_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_4_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_4_Im <= input_delay_registers_0_4_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_4_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_5_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_5_Re <= input_delay_registers_0_5_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_5_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_5_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_5_Im <= input_delay_registers_0_5_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_5_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_6_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_6_Re <= input_delay_registers_0_6_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_6_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_6_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_6_Im <= input_delay_registers_0_6_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_6_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_7_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_7_Re <= input_delay_registers_0_7_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_7_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_7_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_7_Im <= input_delay_registers_0_7_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_7_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_8_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_8_Re <= input_delay_registers_0_8_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_8_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_8_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_8_Im <= input_delay_registers_0_8_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_8_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_9_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_9_Re <= input_delay_registers_0_9_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_9_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_9_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_9_Im <= input_delay_registers_0_9_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_9_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_10_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_10_Re <= input_delay_registers_0_10_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_10_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_10_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_10_Im <= input_delay_registers_0_10_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_10_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_11_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_11_Re <= input_delay_registers_0_11_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_11_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_11_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_11_Im <= input_delay_registers_0_11_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_11_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_0_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_0_Re <= input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_0_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_0_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_0_Im <= input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_0_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_1_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_1_Re <= input_delay_registers_1_1_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_1_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_1_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_1_Im <= input_delay_registers_1_1_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_1_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_2_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_2_Re <= input_delay_registers_1_2_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_2_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_2_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_2_Im <= input_delay_registers_1_2_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_2_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_3_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_3_Re <= input_delay_registers_1_3_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_3_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_3_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_3_Im <= input_delay_registers_1_3_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_3_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_4_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_4_Re <= input_delay_registers_1_4_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_4_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_4_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_4_Im <= input_delay_registers_1_4_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_4_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_5_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_5_Re <= input_delay_registers_1_5_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_5_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_5_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_5_Im <= input_delay_registers_1_5_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_5_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_6_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_6_Re <= input_delay_registers_1_6_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_6_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_6_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_6_Im <= input_delay_registers_1_6_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_6_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_7_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_7_Re <= input_delay_registers_1_7_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_7_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_7_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_7_Im <= input_delay_registers_1_7_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_7_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_8_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_8_Re <= input_delay_registers_1_8_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_8_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_8_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_8_Im <= input_delay_registers_1_8_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_8_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_9_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_9_Re <= input_delay_registers_1_9_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_9_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_9_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_9_Im <= input_delay_registers_1_9_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_9_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_10_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_10_Re <= input_delay_registers_1_10_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_10_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_10_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_10_Im <= input_delay_registers_1_10_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_10_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_11_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_11_Re <= input_delay_registers_1_11_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_11_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_2_11_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_2_11_Im <= input_delay_registers_1_11_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_2_11_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_0_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_0_Re <= input_delay_registers_2_0_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_0_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_0_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_0_Im <= input_delay_registers_2_0_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_0_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_1_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_1_Re <= input_delay_registers_2_1_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_1_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_1_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_1_Im <= input_delay_registers_2_1_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_1_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_2_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_2_Re <= input_delay_registers_2_2_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_2_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_2_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_2_Im <= input_delay_registers_2_2_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_2_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_3_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_3_Re <= input_delay_registers_2_3_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_3_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_3_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_3_Im <= input_delay_registers_2_3_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_3_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_4_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_4_Re <= input_delay_registers_2_4_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_4_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_4_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_4_Im <= input_delay_registers_2_4_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_4_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_5_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_5_Re <= input_delay_registers_2_5_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_5_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_5_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_5_Im <= input_delay_registers_2_5_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_5_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_6_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_6_Re <= input_delay_registers_2_6_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_6_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_6_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_6_Im <= input_delay_registers_2_6_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_6_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_7_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_7_Re <= input_delay_registers_2_7_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_7_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_7_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_7_Im <= input_delay_registers_2_7_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_7_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_8_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_8_Re <= input_delay_registers_2_8_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_8_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_8_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_8_Im <= input_delay_registers_2_8_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_8_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_9_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_9_Re <= input_delay_registers_2_9_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_9_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_9_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_9_Im <= input_delay_registers_2_9_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_9_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_10_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_10_Re <= input_delay_registers_2_10_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_10_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_10_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_10_Im <= input_delay_registers_2_10_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_10_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_11_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_11_Re <= input_delay_registers_2_11_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_11_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_3_11_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_3_11_Im <= input_delay_registers_2_11_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_3_11_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2912:25]
      cnt2 <= 4'h0; // @[FFTDesigns.scala 2912:25]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      if (cnt2 == 4'hb & cnt == 3'h7) begin // @[FFTDesigns.scala 2922:69]
        cnt2 <= 4'h0; // @[FFTDesigns.scala 2923:16]
      end else if (_T_3) begin // @[FFTDesigns.scala 2926:47]
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2928:16]
      end else begin
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2931:16]
      end
    end else begin
      cnt2 <= 4'h0; // @[FFTDesigns.scala 3019:14]
    end
    if (reset) begin // @[FFTDesigns.scala 2913:24]
      cnt <= 3'h0; // @[FFTDesigns.scala 2913:24]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      if (cnt2 == 4'hb & cnt == 3'h7) begin // @[FFTDesigns.scala 2922:69]
        cnt <= 3'h0; // @[FFTDesigns.scala 2924:15]
      end else if (!(_T_3)) begin // @[FFTDesigns.scala 2926:47]
        cnt <= _GEN_0;
      end
    end else begin
      cnt <= 3'h0; // @[FFTDesigns.scala 3018:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  input_delay_registers_0_0_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  input_delay_registers_0_0_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  input_delay_registers_0_1_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  input_delay_registers_0_1_Im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  input_delay_registers_0_2_Re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  input_delay_registers_0_2_Im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  input_delay_registers_0_3_Re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  input_delay_registers_0_3_Im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  input_delay_registers_0_4_Re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  input_delay_registers_0_4_Im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  input_delay_registers_0_5_Re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  input_delay_registers_0_5_Im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  input_delay_registers_0_6_Re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  input_delay_registers_0_6_Im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  input_delay_registers_0_7_Re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  input_delay_registers_0_7_Im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  input_delay_registers_0_8_Re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  input_delay_registers_0_8_Im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  input_delay_registers_0_9_Re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  input_delay_registers_0_9_Im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  input_delay_registers_0_10_Re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  input_delay_registers_0_10_Im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  input_delay_registers_0_11_Re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  input_delay_registers_0_11_Im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  input_delay_registers_1_0_Re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  input_delay_registers_1_0_Im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  input_delay_registers_1_1_Re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  input_delay_registers_1_1_Im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  input_delay_registers_1_2_Re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  input_delay_registers_1_2_Im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  input_delay_registers_1_3_Re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  input_delay_registers_1_3_Im = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  input_delay_registers_1_4_Re = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  input_delay_registers_1_4_Im = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  input_delay_registers_1_5_Re = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  input_delay_registers_1_5_Im = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  input_delay_registers_1_6_Re = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  input_delay_registers_1_6_Im = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  input_delay_registers_1_7_Re = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  input_delay_registers_1_7_Im = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  input_delay_registers_1_8_Re = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  input_delay_registers_1_8_Im = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  input_delay_registers_1_9_Re = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  input_delay_registers_1_9_Im = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  input_delay_registers_1_10_Re = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  input_delay_registers_1_10_Im = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  input_delay_registers_1_11_Re = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  input_delay_registers_1_11_Im = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  input_delay_registers_2_0_Re = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  input_delay_registers_2_0_Im = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  input_delay_registers_2_1_Re = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  input_delay_registers_2_1_Im = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  input_delay_registers_2_2_Re = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  input_delay_registers_2_2_Im = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  input_delay_registers_2_3_Re = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  input_delay_registers_2_3_Im = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  input_delay_registers_2_4_Re = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  input_delay_registers_2_4_Im = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  input_delay_registers_2_5_Re = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  input_delay_registers_2_5_Im = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  input_delay_registers_2_6_Re = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  input_delay_registers_2_6_Im = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  input_delay_registers_2_7_Re = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  input_delay_registers_2_7_Im = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  input_delay_registers_2_8_Re = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  input_delay_registers_2_8_Im = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  input_delay_registers_2_9_Re = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  input_delay_registers_2_9_Im = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  input_delay_registers_2_10_Re = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  input_delay_registers_2_10_Im = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  input_delay_registers_2_11_Re = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  input_delay_registers_2_11_Im = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  input_delay_registers_3_0_Re = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  input_delay_registers_3_0_Im = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  input_delay_registers_3_1_Re = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  input_delay_registers_3_1_Im = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  input_delay_registers_3_2_Re = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  input_delay_registers_3_2_Im = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  input_delay_registers_3_3_Re = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  input_delay_registers_3_3_Im = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  input_delay_registers_3_4_Re = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  input_delay_registers_3_4_Im = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  input_delay_registers_3_5_Re = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  input_delay_registers_3_5_Im = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  input_delay_registers_3_6_Re = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  input_delay_registers_3_6_Im = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  input_delay_registers_3_7_Re = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  input_delay_registers_3_7_Im = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  input_delay_registers_3_8_Re = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  input_delay_registers_3_8_Im = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  input_delay_registers_3_9_Re = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  input_delay_registers_3_9_Im = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  input_delay_registers_3_10_Re = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  input_delay_registers_3_10_Im = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  input_delay_registers_3_11_Re = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  input_delay_registers_3_11_Im = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  cnt2 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  cnt = _RAND_98[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_mr(
  input  [6:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_2_Re,
  output [31:0] io_out_data_2_Im,
  output [31:0] io_out_data_4_Re,
  output [31:0] io_out_data_4_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_8_Re,
  output [31:0] io_out_data_8_Im,
  output [31:0] io_out_data_10_Re,
  output [31:0] io_out_data_10_Im,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_11_Im
);
  wire [31:0] _GEN_17 = 3'h1 == io_in_addr[2:0] ? 32'h3f7746ea : 32'h3f800000; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_18 = 3'h2 == io_in_addr[2:0] ? 32'h3f5db3d6 : _GEN_17; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_19 = 3'h3 == io_in_addr[2:0] ? 32'h3f3504f2 : _GEN_18; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_20 = 3'h4 == io_in_addr[2:0] ? 32'h3f000000 : _GEN_19; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_21 = 3'h5 == io_in_addr[2:0] ? 32'h3e8483ec : _GEN_20; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_22 = 3'h6 == io_in_addr[2:0] ? 32'h248d3131 : _GEN_21; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_25 = 3'h1 == io_in_addr[2:0] ? 32'hbe8483ec : 32'h80800000; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_26 = 3'h2 == io_in_addr[2:0] ? 32'hbefffffc : _GEN_25; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_27 = 3'h3 == io_in_addr[2:0] ? 32'hbf3504f2 : _GEN_26; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_28 = 3'h4 == io_in_addr[2:0] ? 32'hbf5db3d6 : _GEN_27; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_29 = 3'h5 == io_in_addr[2:0] ? 32'hbf7746ea : _GEN_28; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_30 = 3'h6 == io_in_addr[2:0] ? 32'hbf800000 : _GEN_29; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_33 = 3'h1 == io_in_addr[2:0] ? 32'h3f5db3d6 : 32'h3f800000; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_34 = 3'h2 == io_in_addr[2:0] ? 32'h3f000000 : _GEN_33; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_35 = 3'h3 == io_in_addr[2:0] ? 32'h248d3131 : _GEN_34; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_36 = 3'h4 == io_in_addr[2:0] ? 32'hbefffffc : _GEN_35; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_37 = 3'h5 == io_in_addr[2:0] ? 32'hbf5db3d6 : _GEN_36; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_38 = 3'h6 == io_in_addr[2:0] ? 32'hbf800000 : _GEN_37; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_41 = 3'h1 == io_in_addr[2:0] ? 32'hbefffffc : 32'h80800000; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_42 = 3'h2 == io_in_addr[2:0] ? 32'hbf5db3d6 : _GEN_41; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_43 = 3'h3 == io_in_addr[2:0] ? 32'hbf800000 : _GEN_42; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_44 = 3'h4 == io_in_addr[2:0] ? 32'hbf5db3d6 : _GEN_43; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_45 = 3'h5 == io_in_addr[2:0] ? 32'hbf000000 : _GEN_44; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_46 = 3'h6 == io_in_addr[2:0] ? 32'ha50d3131 : _GEN_45; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_65 = 3'h1 == io_in_addr[2:0] ? 32'h3f726a02 : 32'h3f7f73ae; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_66 = 3'h2 == io_in_addr[2:0] ? 32'h3f54db30 : _GEN_65; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_67 = 3'h3 == io_in_addr[2:0] ? 32'h3f28cae2 : _GEN_66; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_68 = 3'h4 == io_in_addr[2:0] ? 32'h3ee273a8 : _GEN_67; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_69 = 3'h5 == io_in_addr[2:0] ? 32'h3e47c5c0 : _GEN_68; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_70 = 3'h6 == io_in_addr[2:0] ? 32'hbd85f210 : _GEN_69; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_73 = 3'h1 == io_in_addr[2:0] ? 32'hbea493b4 : 32'hbd85f210; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_74 = 3'h2 == io_in_addr[2:0] ? 32'hbf0e39d8 : _GEN_73; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_75 = 3'h3 == io_in_addr[2:0] ? 32'hbf407892 : _GEN_74; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_76 = 3'h4 == io_in_addr[2:0] ? 32'hbf659972 : _GEN_75; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_77 = 3'h5 == io_in_addr[2:0] ? 32'hbf7b14be : _GEN_76; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_78 = 3'h6 == io_in_addr[2:0] ? 32'hbf7f73ae : _GEN_77; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_81 = 3'h1 == io_in_addr[2:0] ? 32'h3f4b1934 : 32'h3f7dcf54; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_82 = 3'h2 == io_in_addr[2:0] ? 32'h3ec3ef14 : _GEN_81; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_83 = 3'h3 == io_in_addr[2:0] ? 32'hbe05a8a8 : _GEN_82; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_84 = 3'h4 == io_in_addr[2:0] ? 32'hbf1bd7c8 : _GEN_83; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_85 = 3'h5 == io_in_addr[2:0] ? 32'hbf6c835e : _GEN_84; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_86 = 3'h6 == io_in_addr[2:0] ? 32'hbf7dcf54 : _GEN_85; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_89 = 3'h1 == io_in_addr[2:0] ? 32'hbf1bd7c8 : 32'hbe05a8a8; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_90 = 3'h2 == io_in_addr[2:0] ? 32'hbf6c835e : _GEN_89; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_91 = 3'h3 == io_in_addr[2:0] ? 32'hbf7dcf54 : _GEN_90; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_92 = 3'h4 == io_in_addr[2:0] ? 32'hbf4b1934 : _GEN_91; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_93 = 3'h5 == io_in_addr[2:0] ? 32'hbec3ef14 : _GEN_92; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_94 = 3'h6 == io_in_addr[2:0] ? 32'h3e05a8a8 : _GEN_93; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_113 = 3'h1 == io_in_addr[2:0] ? 32'h3f6c835e : 32'h3f7dcf54; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_114 = 3'h2 == io_in_addr[2:0] ? 32'h3f4b1934 : _GEN_113; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_115 = 3'h3 == io_in_addr[2:0] ? 32'h3f1bd7c8 : _GEN_114; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_116 = 3'h4 == io_in_addr[2:0] ? 32'h3ec3ef14 : _GEN_115; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_117 = 3'h5 == io_in_addr[2:0] ? 32'h3e05a8a8 : _GEN_116; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_118 = 3'h6 == io_in_addr[2:0] ? 32'hbe05a8a8 : _GEN_117; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_121 = 3'h1 == io_in_addr[2:0] ? 32'hbec3ef14 : 32'hbe05a8a8; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_122 = 3'h2 == io_in_addr[2:0] ? 32'hbf1bd7c8 : _GEN_121; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_123 = 3'h3 == io_in_addr[2:0] ? 32'hbf4b1934 : _GEN_122; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_124 = 3'h4 == io_in_addr[2:0] ? 32'hbf6c835e : _GEN_123; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_125 = 3'h5 == io_in_addr[2:0] ? 32'hbf7dcf54 : _GEN_124; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_126 = 3'h6 == io_in_addr[2:0] ? 32'hbf7dcf54 : _GEN_125; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_129 = 3'h1 == io_in_addr[2:0] ? 32'h3f3504f2 : 32'h3f7746ea; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_130 = 3'h2 == io_in_addr[2:0] ? 32'h3e8483ec : _GEN_129; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_131 = 3'h3 == io_in_addr[2:0] ? 32'hbe8483ec : _GEN_130; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_132 = 3'h4 == io_in_addr[2:0] ? 32'hbf3504f2 : _GEN_131; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_133 = 3'h5 == io_in_addr[2:0] ? 32'hbf7746ea : _GEN_132; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_134 = 3'h6 == io_in_addr[2:0] ? 32'hbf7746ea : _GEN_133; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_137 = 3'h1 == io_in_addr[2:0] ? 32'hbf3504f2 : 32'hbe8483ec; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_138 = 3'h2 == io_in_addr[2:0] ? 32'hbf7746ea : _GEN_137; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_139 = 3'h3 == io_in_addr[2:0] ? 32'hbf7746ea : _GEN_138; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_140 = 3'h4 == io_in_addr[2:0] ? 32'hbf3504f2 : _GEN_139; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_141 = 3'h5 == io_in_addr[2:0] ? 32'hbe8483ec : _GEN_140; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_142 = 3'h6 == io_in_addr[2:0] ? 32'h3e8483ec : _GEN_141; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_161 = 3'h1 == io_in_addr[2:0] ? 32'h3f659972 : 32'h3f7b14be; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_162 = 3'h2 == io_in_addr[2:0] ? 32'h3f407892 : _GEN_161; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_163 = 3'h3 == io_in_addr[2:0] ? 32'h3f0e39d8 : _GEN_162; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_164 = 3'h4 == io_in_addr[2:0] ? 32'h3ea493b4 : _GEN_163; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_165 = 3'h5 == io_in_addr[2:0] ? 32'h3d85f210 : _GEN_164; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_166 = 3'h6 == io_in_addr[2:0] ? 32'hbe47c5c0 : _GEN_165; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_169 = 3'h1 == io_in_addr[2:0] ? 32'hbee273a8 : 32'hbe47c5c0; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_170 = 3'h2 == io_in_addr[2:0] ? 32'hbf28cae2 : _GEN_169; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_171 = 3'h3 == io_in_addr[2:0] ? 32'hbf54db30 : _GEN_170; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_172 = 3'h4 == io_in_addr[2:0] ? 32'hbf726a02 : _GEN_171; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_173 = 3'h5 == io_in_addr[2:0] ? 32'hbf7f73ae : _GEN_172; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_174 = 3'h6 == io_in_addr[2:0] ? 32'hbf7b14be : _GEN_173; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_177 = 3'h1 == io_in_addr[2:0] ? 32'h3f1bd7c8 : 32'h3f6c835e; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_178 = 3'h2 == io_in_addr[2:0] ? 32'h3e05a8a8 : _GEN_177; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_179 = 3'h3 == io_in_addr[2:0] ? 32'hbec3ef14 : _GEN_178; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_180 = 3'h4 == io_in_addr[2:0] ? 32'hbf4b1934 : _GEN_179; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_181 = 3'h5 == io_in_addr[2:0] ? 32'hbf7dcf54 : _GEN_180; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_182 = 3'h6 == io_in_addr[2:0] ? 32'hbf6c835e : _GEN_181; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_185 = 3'h1 == io_in_addr[2:0] ? 32'hbf4b1934 : 32'hbec3ef14; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_186 = 3'h2 == io_in_addr[2:0] ? 32'hbf7dcf54 : _GEN_185; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_187 = 3'h3 == io_in_addr[2:0] ? 32'hbf6c835e : _GEN_186; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_188 = 3'h4 == io_in_addr[2:0] ? 32'hbf1bd7c8 : _GEN_187; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_189 = 3'h5 == io_in_addr[2:0] ? 32'hbe05a8a8 : _GEN_188; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_190 = 3'h6 == io_in_addr[2:0] ? 32'h3ec3ef14 : _GEN_189; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_1_Re = 3'h7 == io_in_addr[2:0] ? 32'hbe8483ec : _GEN_22; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_1_Im = 3'h7 == io_in_addr[2:0] ? 32'hbf7746ea : _GEN_30; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_2_Re = 3'h7 == io_in_addr[2:0] ? 32'hbf5db3d6 : _GEN_38; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_2_Im = 3'h7 == io_in_addr[2:0] ? 32'h3efffffc : _GEN_46; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_4_Re = 3'h7 == io_in_addr[2:0] ? 32'hbea493b4 : _GEN_70; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_4_Im = 3'h7 == io_in_addr[2:0] ? 32'hbf726a02 : _GEN_78; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_5_Re = 3'h7 == io_in_addr[2:0] ? 32'hbf4b1934 : _GEN_86; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_5_Im = 3'h7 == io_in_addr[2:0] ? 32'h3f1bd7c8 : _GEN_94; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_7_Re = 3'h7 == io_in_addr[2:0] ? 32'hbec3ef14 : _GEN_118; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_7_Im = 3'h7 == io_in_addr[2:0] ? 32'hbf6c835e : _GEN_126; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_8_Re = 3'h7 == io_in_addr[2:0] ? 32'hbf3504f2 : _GEN_134; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_8_Im = 3'h7 == io_in_addr[2:0] ? 32'h3f3504f2 : _GEN_142; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_10_Re = 3'h7 == io_in_addr[2:0] ? 32'hbee273a8 : _GEN_166; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_10_Im = 3'h7 == io_in_addr[2:0] ? 32'hbf659972 : _GEN_174; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_11_Re = 3'h7 == io_in_addr[2:0] ? 32'hbf1bd7c8 : _GEN_182; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_11_Im = 3'h7 == io_in_addr[2:0] ? 32'h3f4b1934 : _GEN_190; // @[FFTDesigns.scala 2085:{25,25}]
endmodule
module TwiddleFactorsStreamed_mr_v2(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] TwiddleFactorROM_mr_io_in_addr; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_1_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_1_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_2_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_2_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_4_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_4_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_5_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_5_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_7_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_7_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_8_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_8_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_10_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_10_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_11_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_11_Im; // @[FFTDesigns.scala 2314:26]
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_1_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_2_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_3_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_4_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_5_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_6_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_7_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_8_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_8_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_9_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_9_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_10_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_10_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_11_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_11_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  reg [2:0] cnt; // @[FFTDesigns.scala 2322:24]
  reg [3:0] cnt2; // @[FFTDesigns.scala 2323:25]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2324:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2324:28]
  wire [3:0] _cnt2_T_1 = cnt2 + 4'h1; // @[FFTDesigns.scala 2339:24]
  wire [2:0] _cnt_T_1 = cnt + 3'h1; // @[FFTDesigns.scala 2341:22]
  TwiddleFactorROM_mr TwiddleFactorROM_mr ( // @[FFTDesigns.scala 2314:26]
    .io_in_addr(TwiddleFactorROM_mr_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_mr_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_mr_io_out_data_1_Im),
    .io_out_data_2_Re(TwiddleFactorROM_mr_io_out_data_2_Re),
    .io_out_data_2_Im(TwiddleFactorROM_mr_io_out_data_2_Im),
    .io_out_data_4_Re(TwiddleFactorROM_mr_io_out_data_4_Re),
    .io_out_data_4_Im(TwiddleFactorROM_mr_io_out_data_4_Im),
    .io_out_data_5_Re(TwiddleFactorROM_mr_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_mr_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_mr_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_mr_io_out_data_7_Im),
    .io_out_data_8_Re(TwiddleFactorROM_mr_io_out_data_8_Re),
    .io_out_data_8_Im(TwiddleFactorROM_mr_io_out_data_8_Im),
    .io_out_data_10_Re(TwiddleFactorROM_mr_io_out_data_10_Re),
    .io_out_data_10_Im(TwiddleFactorROM_mr_io_out_data_10_Im),
    .io_out_data_11_Re(TwiddleFactorROM_mr_io_out_data_11_Re),
    .io_out_data_11_Im(TwiddleFactorROM_mr_io_out_data_11_Im)
  );
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_clock),
    .reset(FPComplexMult_reset),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_1_clock),
    .reset(FPComplexMult_1_reset),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_2_clock),
    .reset(FPComplexMult_2_reset),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_3_clock),
    .reset(FPComplexMult_3_reset),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_4_clock),
    .reset(FPComplexMult_4_reset),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_5_clock),
    .reset(FPComplexMult_5_reset),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_6_clock),
    .reset(FPComplexMult_6_reset),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_7_clock),
    .reset(FPComplexMult_7_reset),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_8 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_8_clock),
    .reset(FPComplexMult_8_reset),
    .io_in_a_Re(FPComplexMult_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_8_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_9 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_9_clock),
    .reset(FPComplexMult_9_reset),
    .io_in_a_Re(FPComplexMult_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_9_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_10 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_10_clock),
    .reset(FPComplexMult_10_reset),
    .io_in_a_Re(FPComplexMult_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_10_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_11 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_11_clock),
    .reset(FPComplexMult_11_reset),
    .io_in_a_Re(FPComplexMult_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_11_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_8_Re = FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_8_Im = FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_9_Re = FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_9_Im = FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_10_Re = FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_10_Im = FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_11_Re = FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_11_Im = FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign TwiddleFactorROM_mr_io_in_addr = {{4'd0}, cnt}; // @[FFTDesigns.scala 2359:24]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_reset = reset;
  assign FPComplexMult_io_in_a_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_io_in_a_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_reset = reset;
  assign FPComplexMult_1_io_in_a_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_1_io_in_a_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_1_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_1_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_1_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_1_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_reset = reset;
  assign FPComplexMult_2_io_in_a_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_2_io_in_a_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_2_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_2_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_2_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_2_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_reset = reset;
  assign FPComplexMult_3_io_in_a_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_3_io_in_a_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_3_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_3_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_reset = reset;
  assign FPComplexMult_4_io_in_a_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_4_io_in_a_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_4_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_4_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_4_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_4_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_reset = reset;
  assign FPComplexMult_5_io_in_a_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_5_io_in_a_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_5_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_5_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_5_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_5_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_reset = reset;
  assign FPComplexMult_6_io_in_a_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_6_io_in_a_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_6_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_6_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_reset = reset;
  assign FPComplexMult_7_io_in_a_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_7_io_in_a_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_7_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_7_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_7_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_7_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_8_clock = clock;
  assign FPComplexMult_8_reset = reset;
  assign FPComplexMult_8_io_in_a_Re = _T_1 ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_8_io_in_a_Im = _T_1 ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_8_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_8_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_8_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_8_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_9_clock = clock;
  assign FPComplexMult_9_reset = reset;
  assign FPComplexMult_9_io_in_a_Re = _T_1 ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_9_io_in_a_Im = _T_1 ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_9_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_9_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_10_clock = clock;
  assign FPComplexMult_10_reset = reset;
  assign FPComplexMult_10_io_in_a_Re = _T_1 ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_10_io_in_a_Im = _T_1 ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_10_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_10_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_10_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_10_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_11_clock = clock;
  assign FPComplexMult_11_reset = reset;
  assign FPComplexMult_11_io_in_a_Re = _T_1 ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_11_io_in_a_Im = _T_1 ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_11_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_11_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_11_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_11_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2322:24]
      cnt <= 3'h0; // @[FFTDesigns.scala 2322:24]
    end else if (_T_1) begin // @[FFTDesigns.scala 2333:32]
      if (cnt2 == 4'hb) begin // @[FFTDesigns.scala 2334:37]
        cnt <= 3'h0; // @[FFTDesigns.scala 2336:15]
      end else if (!(cnt == 3'h7 & cnt2 != 4'hb)) begin // @[FFTDesigns.scala 2337:66]
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2341:15]
      end
    end else begin
      cnt <= 3'h0; // @[FFTDesigns.scala 2353:13]
    end
    if (reset) begin // @[FFTDesigns.scala 2323:25]
      cnt2 <= 4'h0; // @[FFTDesigns.scala 2323:25]
    end else if (_T_1) begin // @[FFTDesigns.scala 2333:32]
      if (cnt2 == 4'hb) begin // @[FFTDesigns.scala 2334:37]
        cnt2 <= 4'h0; // @[FFTDesigns.scala 2335:16]
      end else if (cnt == 3'h7 & cnt2 != 4'hb) begin // @[FFTDesigns.scala 2337:66]
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2339:16]
      end else begin
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2342:16]
      end
    end else begin
      cnt2 <= 4'h0; // @[FFTDesigns.scala 2354:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  cnt2 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module od_fft96_8_12(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input         io_in_ready,
  output        io_out_validate,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
`endif // RANDOMIZE_REG_INIT
  wire  FFT_sr_v2_streaming_nrv_clock; // @[FFTDesigns.scala 6453:32]
  wire  FFT_sr_v2_streaming_nrv_reset; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_0_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_0_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_1_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_1_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_2_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_2_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_3_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_3_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_4_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_4_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_5_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_5_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_6_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_6_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_7_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_7_Im; // @[FFTDesigns.scala 6453:32]
  wire  FFT_sr_v2_streaming_nrv_io_in_ready; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_0_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_0_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_1_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_1_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_2_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_2_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_3_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_3_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_4_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_4_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_5_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_5_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_6_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_6_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_7_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_7_Im; // @[FFTDesigns.scala 6453:32]
  wire  DFT_r_v2_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_1_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_1_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_2_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_2_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_3_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_3_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  PermutationsWithStreaming_clock; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_reset; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_0_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_0_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_1_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_1_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_2_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_2_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_3_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_3_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_4_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_4_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_5_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_5_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_6_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_6_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_7_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_7_Im; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_0; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_1; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_2; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_3; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_4; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_5; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_6; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_7; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_8; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_9; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_10; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_11; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_12; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_13; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_14; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_15; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_16; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_17; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_18; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_19; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_20; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_21; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_22; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_23; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_24; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_0_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_0_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_1_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_1_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_2_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_2_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_3_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_3_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_4_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_4_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_5_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_5_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_6_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_6_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_7_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_7_Im; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_mr_clock; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_reset; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_0_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_0_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_1_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_1_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_2_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_2_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_3_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_3_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_4_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_4_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_5_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_5_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_6_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_6_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_7_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_7_Im; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_0; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_1; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_2; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_3; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_4; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_5; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_6; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_7; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_8; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_9; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_10; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_11; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_12; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_13; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_14; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_15; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_16; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_17; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_18; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_19; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_20; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_21; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_22; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_23; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_24; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_0_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_0_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_1_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_1_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_2_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_2_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_3_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_3_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_4_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_4_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_5_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_5_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_6_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_6_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_7_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_7_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_8_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_8_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_9_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_9_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_10_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_10_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_11_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_11_Im; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_1_clock; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_reset; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_0_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_0_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_1_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_1_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_2_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_2_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_3_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_3_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_4_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_4_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_5_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_5_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_6_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_6_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_7_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_7_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_8_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_8_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_9_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_9_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_10_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_10_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_11_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_11_Im; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_0; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_1; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_2; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_3; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_4; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_5; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_6; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_7; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_8; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_9; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_10; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_11; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_12; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_13; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_14; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_15; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_16; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_17; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_18; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_19; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_20; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_21; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_22; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_23; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_24; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_0_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_0_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_1_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_1_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_2_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_2_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_3_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_3_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_4_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_4_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_5_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_5_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_6_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_6_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_7_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_7_Im; // @[FFTDesigns.scala 6470:32]
  wire  TwiddleFactorsStreamed_mr_v2_clock; // @[FFTDesigns.scala 6471:32]
  wire  TwiddleFactorsStreamed_mr_v2_reset; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_0_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_0_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_1_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_1_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_2_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_2_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_3_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_3_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_4_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_4_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_5_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_5_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_6_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_6_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_7_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_7_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_8_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_8_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_9_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_9_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_10_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_10_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_11_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_11_Im; // @[FFTDesigns.scala 6471:32]
  wire  TwiddleFactorsStreamed_mr_v2_io_in_en_0; // @[FFTDesigns.scala 6471:32]
  wire  TwiddleFactorsStreamed_mr_v2_io_in_en_1; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_0_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_0_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_1_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_1_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_2_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_2_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_3_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_3_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_4_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_4_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_5_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_5_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_6_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_6_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_7_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_7_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_8_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_8_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_9_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_9_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_10_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_10_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_11_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_11_Im; // @[FFTDesigns.scala 6471:32]
  reg  DFT_regdelays1_0; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_1; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_2; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_3; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_4; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_5; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_6; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_7; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_8; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_9; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_10; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_11; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_12; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_13; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_14; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_15; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_16; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_17; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_18; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_19; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_20; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_21; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_22; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_23; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_24; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_25; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_26; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_27; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_28; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_29; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_30; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_31; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_32; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_33; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_34; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_35; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_36; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_37; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_38; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_39; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_40; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_41; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_42; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_43; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_44; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_45; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_46; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_47; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_48; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_49; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_50; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_51; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_52; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_53; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_54; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_55; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_56; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_57; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_58; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_59; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_60; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays2_0; // @[FFTDesigns.scala 6475:35]
  reg  DFT_regdelays2_1; // @[FFTDesigns.scala 6475:35]
  reg  DFT_regdelays2_2; // @[FFTDesigns.scala 6475:35]
  reg  DFT_regdelays2_3; // @[FFTDesigns.scala 6475:35]
  reg  Twid_regdelays_0; // @[FFTDesigns.scala 6476:35]
  reg  Twid_regdelays_1; // @[FFTDesigns.scala 6476:35]
  reg  Perm_regdelays1_0_0; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_1; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_2; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_3; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_4; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_5; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_6; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_7; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_8; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_9; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_10; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_11; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_12; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_13; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_14; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_15; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_16; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_17; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_18; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_19; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_20; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_21; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_22; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_23; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_0; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_1; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_2; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_3; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_4; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_5; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_6; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_7; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_8; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_9; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_10; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_11; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_12; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_13; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_14; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_15; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_16; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_17; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_18; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_19; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_20; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_21; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_22; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_23; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_0; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_1; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_2; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_3; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_4; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_5; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_6; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_7; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_8; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_9; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_10; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_11; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_12; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_13; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_14; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_15; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_16; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_17; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_18; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_19; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_20; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_21; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_22; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_23; // @[FFTDesigns.scala 6477:36]
  reg  out_regdelay; // @[FFTDesigns.scala 6478:33]
  reg [31:0] results_0_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_0_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_1_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_1_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_2_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_2_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_3_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_3_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_4_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_4_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_5_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_5_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_6_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_6_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_7_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_7_Im; // @[FFTDesigns.scala 6479:28]
  FFT_sr_v2_streaming_nrv FFT_sr_v2_streaming_nrv ( // @[FFTDesigns.scala 6453:32]
    .clock(FFT_sr_v2_streaming_nrv_clock),
    .reset(FFT_sr_v2_streaming_nrv_reset),
    .io_in_0_Re(FFT_sr_v2_streaming_nrv_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_streaming_nrv_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_streaming_nrv_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_streaming_nrv_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_streaming_nrv_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_streaming_nrv_io_in_2_Im),
    .io_in_3_Re(FFT_sr_v2_streaming_nrv_io_in_3_Re),
    .io_in_3_Im(FFT_sr_v2_streaming_nrv_io_in_3_Im),
    .io_in_4_Re(FFT_sr_v2_streaming_nrv_io_in_4_Re),
    .io_in_4_Im(FFT_sr_v2_streaming_nrv_io_in_4_Im),
    .io_in_5_Re(FFT_sr_v2_streaming_nrv_io_in_5_Re),
    .io_in_5_Im(FFT_sr_v2_streaming_nrv_io_in_5_Im),
    .io_in_6_Re(FFT_sr_v2_streaming_nrv_io_in_6_Re),
    .io_in_6_Im(FFT_sr_v2_streaming_nrv_io_in_6_Im),
    .io_in_7_Re(FFT_sr_v2_streaming_nrv_io_in_7_Re),
    .io_in_7_Im(FFT_sr_v2_streaming_nrv_io_in_7_Im),
    .io_in_ready(FFT_sr_v2_streaming_nrv_io_in_ready),
    .io_out_0_Re(FFT_sr_v2_streaming_nrv_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_streaming_nrv_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_streaming_nrv_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_streaming_nrv_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_streaming_nrv_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_streaming_nrv_io_out_2_Im),
    .io_out_3_Re(FFT_sr_v2_streaming_nrv_io_out_3_Re),
    .io_out_3_Im(FFT_sr_v2_streaming_nrv_io_out_3_Im),
    .io_out_4_Re(FFT_sr_v2_streaming_nrv_io_out_4_Re),
    .io_out_4_Im(FFT_sr_v2_streaming_nrv_io_out_4_Im),
    .io_out_5_Re(FFT_sr_v2_streaming_nrv_io_out_5_Re),
    .io_out_5_Im(FFT_sr_v2_streaming_nrv_io_out_5_Im),
    .io_out_6_Re(FFT_sr_v2_streaming_nrv_io_out_6_Re),
    .io_out_6_Im(FFT_sr_v2_streaming_nrv_io_out_6_Im),
    .io_out_7_Re(FFT_sr_v2_streaming_nrv_io_out_7_Re),
    .io_out_7_Im(FFT_sr_v2_streaming_nrv_io_out_7_Im)
  );
  DFT_r_v2_20 DFT_r_v2 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_clock),
    .reset(DFT_r_v2_reset),
    .io_in_0_Re(DFT_r_v2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_io_out_2_Im)
  );
  DFT_r_v2_20 DFT_r_v2_1 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_1_clock),
    .reset(DFT_r_v2_1_reset),
    .io_in_0_Re(DFT_r_v2_1_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_1_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_1_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_1_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_1_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_1_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_1_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_1_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_1_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_1_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_1_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_1_io_out_2_Im)
  );
  DFT_r_v2_20 DFT_r_v2_2 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_2_clock),
    .reset(DFT_r_v2_2_reset),
    .io_in_0_Re(DFT_r_v2_2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_2_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_2_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_2_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_2_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_2_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_2_io_out_2_Im)
  );
  DFT_r_v2_20 DFT_r_v2_3 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_3_clock),
    .reset(DFT_r_v2_3_reset),
    .io_in_0_Re(DFT_r_v2_3_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_3_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_3_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_3_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_3_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_3_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_3_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_3_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_3_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_3_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_3_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_3_io_out_2_Im)
  );
  PermutationsWithStreaming_6 PermutationsWithStreaming ( // @[FFTDesigns.scala 6468:32]
    .clock(PermutationsWithStreaming_clock),
    .reset(PermutationsWithStreaming_reset),
    .io_in_0_Re(PermutationsWithStreaming_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_io_in_7_Im),
    .io_in_en_0(PermutationsWithStreaming_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_io_in_en_8),
    .io_in_en_9(PermutationsWithStreaming_io_in_en_9),
    .io_in_en_10(PermutationsWithStreaming_io_in_en_10),
    .io_in_en_11(PermutationsWithStreaming_io_in_en_11),
    .io_in_en_12(PermutationsWithStreaming_io_in_en_12),
    .io_in_en_13(PermutationsWithStreaming_io_in_en_13),
    .io_in_en_14(PermutationsWithStreaming_io_in_en_14),
    .io_in_en_15(PermutationsWithStreaming_io_in_en_15),
    .io_in_en_16(PermutationsWithStreaming_io_in_en_16),
    .io_in_en_17(PermutationsWithStreaming_io_in_en_17),
    .io_in_en_18(PermutationsWithStreaming_io_in_en_18),
    .io_in_en_19(PermutationsWithStreaming_io_in_en_19),
    .io_in_en_20(PermutationsWithStreaming_io_in_en_20),
    .io_in_en_21(PermutationsWithStreaming_io_in_en_21),
    .io_in_en_22(PermutationsWithStreaming_io_in_en_22),
    .io_in_en_23(PermutationsWithStreaming_io_in_en_23),
    .io_in_en_24(PermutationsWithStreaming_io_in_en_24),
    .io_out_0_Re(PermutationsWithStreaming_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_io_out_7_Im)
  );
  PermutationsWithStreaming_mr PermutationsWithStreaming_mr ( // @[FFTDesigns.scala 6469:32]
    .clock(PermutationsWithStreaming_mr_clock),
    .reset(PermutationsWithStreaming_mr_reset),
    .io_in_0_Re(PermutationsWithStreaming_mr_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_mr_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_mr_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_mr_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_mr_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_mr_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_mr_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_mr_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_mr_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_mr_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_mr_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_mr_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_mr_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_mr_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_mr_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_mr_io_in_7_Im),
    .io_in_en_0(PermutationsWithStreaming_mr_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_mr_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_mr_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_mr_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_mr_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_mr_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_mr_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_mr_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_mr_io_in_en_8),
    .io_in_en_9(PermutationsWithStreaming_mr_io_in_en_9),
    .io_in_en_10(PermutationsWithStreaming_mr_io_in_en_10),
    .io_in_en_11(PermutationsWithStreaming_mr_io_in_en_11),
    .io_in_en_12(PermutationsWithStreaming_mr_io_in_en_12),
    .io_in_en_13(PermutationsWithStreaming_mr_io_in_en_13),
    .io_in_en_14(PermutationsWithStreaming_mr_io_in_en_14),
    .io_in_en_15(PermutationsWithStreaming_mr_io_in_en_15),
    .io_in_en_16(PermutationsWithStreaming_mr_io_in_en_16),
    .io_in_en_17(PermutationsWithStreaming_mr_io_in_en_17),
    .io_in_en_18(PermutationsWithStreaming_mr_io_in_en_18),
    .io_in_en_19(PermutationsWithStreaming_mr_io_in_en_19),
    .io_in_en_20(PermutationsWithStreaming_mr_io_in_en_20),
    .io_in_en_21(PermutationsWithStreaming_mr_io_in_en_21),
    .io_in_en_22(PermutationsWithStreaming_mr_io_in_en_22),
    .io_in_en_23(PermutationsWithStreaming_mr_io_in_en_23),
    .io_in_en_24(PermutationsWithStreaming_mr_io_in_en_24),
    .io_out_0_Re(PermutationsWithStreaming_mr_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_mr_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_mr_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_mr_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_mr_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_mr_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_mr_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_mr_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_mr_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_mr_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_mr_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_mr_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_mr_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_mr_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_mr_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_mr_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_mr_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_mr_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_mr_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_mr_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_mr_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_mr_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_mr_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_mr_io_out_11_Im)
  );
  PermutationsWithStreaming_mr_1 PermutationsWithStreaming_mr_1 ( // @[FFTDesigns.scala 6470:32]
    .clock(PermutationsWithStreaming_mr_1_clock),
    .reset(PermutationsWithStreaming_mr_1_reset),
    .io_in_0_Re(PermutationsWithStreaming_mr_1_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_mr_1_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_mr_1_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_mr_1_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_mr_1_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_mr_1_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_mr_1_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_mr_1_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_mr_1_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_mr_1_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_mr_1_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_mr_1_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_mr_1_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_mr_1_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_mr_1_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_mr_1_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_mr_1_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_mr_1_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_mr_1_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_mr_1_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_mr_1_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_mr_1_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_mr_1_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_mr_1_io_in_11_Im),
    .io_in_en_0(PermutationsWithStreaming_mr_1_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_mr_1_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_mr_1_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_mr_1_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_mr_1_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_mr_1_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_mr_1_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_mr_1_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_mr_1_io_in_en_8),
    .io_in_en_9(PermutationsWithStreaming_mr_1_io_in_en_9),
    .io_in_en_10(PermutationsWithStreaming_mr_1_io_in_en_10),
    .io_in_en_11(PermutationsWithStreaming_mr_1_io_in_en_11),
    .io_in_en_12(PermutationsWithStreaming_mr_1_io_in_en_12),
    .io_in_en_13(PermutationsWithStreaming_mr_1_io_in_en_13),
    .io_in_en_14(PermutationsWithStreaming_mr_1_io_in_en_14),
    .io_in_en_15(PermutationsWithStreaming_mr_1_io_in_en_15),
    .io_in_en_16(PermutationsWithStreaming_mr_1_io_in_en_16),
    .io_in_en_17(PermutationsWithStreaming_mr_1_io_in_en_17),
    .io_in_en_18(PermutationsWithStreaming_mr_1_io_in_en_18),
    .io_in_en_19(PermutationsWithStreaming_mr_1_io_in_en_19),
    .io_in_en_20(PermutationsWithStreaming_mr_1_io_in_en_20),
    .io_in_en_21(PermutationsWithStreaming_mr_1_io_in_en_21),
    .io_in_en_22(PermutationsWithStreaming_mr_1_io_in_en_22),
    .io_in_en_23(PermutationsWithStreaming_mr_1_io_in_en_23),
    .io_in_en_24(PermutationsWithStreaming_mr_1_io_in_en_24),
    .io_out_0_Re(PermutationsWithStreaming_mr_1_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_mr_1_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_mr_1_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_mr_1_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_mr_1_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_mr_1_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_mr_1_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_mr_1_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_mr_1_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_mr_1_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_mr_1_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_mr_1_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_mr_1_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_mr_1_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_mr_1_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_mr_1_io_out_7_Im)
  );
  TwiddleFactorsStreamed_mr_v2 TwiddleFactorsStreamed_mr_v2 ( // @[FFTDesigns.scala 6471:32]
    .clock(TwiddleFactorsStreamed_mr_v2_clock),
    .reset(TwiddleFactorsStreamed_mr_v2_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_mr_v2_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_mr_v2_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_mr_v2_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_mr_v2_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_mr_v2_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_mr_v2_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_mr_v2_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_mr_v2_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_mr_v2_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_mr_v2_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_mr_v2_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_mr_v2_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_mr_v2_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_mr_v2_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_mr_v2_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_mr_v2_io_in_7_Im),
    .io_in_8_Re(TwiddleFactorsStreamed_mr_v2_io_in_8_Re),
    .io_in_8_Im(TwiddleFactorsStreamed_mr_v2_io_in_8_Im),
    .io_in_9_Re(TwiddleFactorsStreamed_mr_v2_io_in_9_Re),
    .io_in_9_Im(TwiddleFactorsStreamed_mr_v2_io_in_9_Im),
    .io_in_10_Re(TwiddleFactorsStreamed_mr_v2_io_in_10_Re),
    .io_in_10_Im(TwiddleFactorsStreamed_mr_v2_io_in_10_Im),
    .io_in_11_Re(TwiddleFactorsStreamed_mr_v2_io_in_11_Re),
    .io_in_11_Im(TwiddleFactorsStreamed_mr_v2_io_in_11_Im),
    .io_in_en_0(TwiddleFactorsStreamed_mr_v2_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_mr_v2_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_mr_v2_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_mr_v2_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_mr_v2_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_mr_v2_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_mr_v2_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_mr_v2_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_mr_v2_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_mr_v2_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_mr_v2_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_mr_v2_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_mr_v2_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_mr_v2_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_mr_v2_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_mr_v2_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_mr_v2_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_mr_v2_io_out_7_Im),
    .io_out_8_Re(TwiddleFactorsStreamed_mr_v2_io_out_8_Re),
    .io_out_8_Im(TwiddleFactorsStreamed_mr_v2_io_out_8_Im),
    .io_out_9_Re(TwiddleFactorsStreamed_mr_v2_io_out_9_Re),
    .io_out_9_Im(TwiddleFactorsStreamed_mr_v2_io_out_9_Im),
    .io_out_10_Re(TwiddleFactorsStreamed_mr_v2_io_out_10_Re),
    .io_out_10_Im(TwiddleFactorsStreamed_mr_v2_io_out_10_Im),
    .io_out_11_Re(TwiddleFactorsStreamed_mr_v2_io_out_11_Re),
    .io_out_11_Im(TwiddleFactorsStreamed_mr_v2_io_out_11_Im)
  );
  assign io_out_validate = out_regdelay; // @[FFTDesigns.scala 6560:23]
  assign io_out_0_Re = results_0_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_0_Im = results_0_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_1_Re = results_1_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_1_Im = results_1_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_2_Re = results_2_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_2_Im = results_2_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_3_Re = results_3_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_3_Im = results_3_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_4_Re = results_4_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_4_Im = results_4_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_5_Re = results_5_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_5_Im = results_5_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_6_Re = results_6_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_6_Im = results_6_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_7_Re = results_7_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_7_Im = results_7_Im; // @[FFTDesigns.scala 6561:14]
  assign FFT_sr_v2_streaming_nrv_clock = clock;
  assign FFT_sr_v2_streaming_nrv_reset = reset;
  assign FFT_sr_v2_streaming_nrv_io_in_0_Re = PermutationsWithStreaming_io_out_0_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_0_Im = PermutationsWithStreaming_io_out_0_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_1_Re = PermutationsWithStreaming_io_out_1_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_1_Im = PermutationsWithStreaming_io_out_1_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_2_Re = PermutationsWithStreaming_io_out_2_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_2_Im = PermutationsWithStreaming_io_out_2_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_3_Re = PermutationsWithStreaming_io_out_3_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_3_Im = PermutationsWithStreaming_io_out_3_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_4_Re = PermutationsWithStreaming_io_out_4_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_4_Im = PermutationsWithStreaming_io_out_4_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_5_Re = PermutationsWithStreaming_io_out_5_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_5_Im = PermutationsWithStreaming_io_out_5_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_6_Re = PermutationsWithStreaming_io_out_6_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_6_Im = PermutationsWithStreaming_io_out_6_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_7_Re = PermutationsWithStreaming_io_out_7_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_7_Im = PermutationsWithStreaming_io_out_7_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_ready = Perm_regdelays1_0_23; // @[FFTDesigns.scala 6536:33]
  assign DFT_r_v2_clock = clock;
  assign DFT_r_v2_reset = reset;
  assign DFT_r_v2_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_0_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_0_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_1_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_1_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_2_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_2_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_clock = clock;
  assign DFT_r_v2_1_reset = reset;
  assign DFT_r_v2_1_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_3_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_3_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_4_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_4_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_5_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_5_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_clock = clock;
  assign DFT_r_v2_2_reset = reset;
  assign DFT_r_v2_2_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_6_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_6_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_7_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_7_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_8_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_8_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_clock = clock;
  assign DFT_r_v2_3_reset = reset;
  assign DFT_r_v2_3_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_9_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_9_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_10_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_10_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_11_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_11_Im; // @[FFTDesigns.scala 6547:37]
  assign PermutationsWithStreaming_clock = clock;
  assign PermutationsWithStreaming_reset = reset;
  assign PermutationsWithStreaming_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_2_Re = io_in_2_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_2_Im = io_in_2_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_3_Re = io_in_3_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_3_Im = io_in_3_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_4_Re = io_in_4_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_4_Im = io_in_4_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_5_Re = io_in_5_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_5_Im = io_in_5_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_6_Re = io_in_6_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_6_Im = io_in_6_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_7_Re = io_in_7_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_7_Im = io_in_7_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_en_0 = io_in_ready; // @[FFTDesigns.scala 6485:37]
  assign PermutationsWithStreaming_io_in_en_1 = Perm_regdelays1_0_0; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_2 = Perm_regdelays1_0_1; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_3 = Perm_regdelays1_0_2; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_4 = Perm_regdelays1_0_3; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_5 = Perm_regdelays1_0_4; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_6 = Perm_regdelays1_0_5; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_7 = Perm_regdelays1_0_6; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_8 = Perm_regdelays1_0_7; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_9 = Perm_regdelays1_0_8; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_10 = Perm_regdelays1_0_9; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_11 = Perm_regdelays1_0_10; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_12 = Perm_regdelays1_0_11; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_13 = Perm_regdelays1_0_12; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_14 = Perm_regdelays1_0_13; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_15 = Perm_regdelays1_0_14; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_16 = Perm_regdelays1_0_15; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_17 = Perm_regdelays1_0_16; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_18 = Perm_regdelays1_0_17; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_19 = Perm_regdelays1_0_18; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_20 = Perm_regdelays1_0_19; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_21 = Perm_regdelays1_0_20; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_22 = Perm_regdelays1_0_21; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_23 = Perm_regdelays1_0_22; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_24 = Perm_regdelays1_0_23; // @[FFTDesigns.scala 6511:51]
  assign PermutationsWithStreaming_mr_clock = clock;
  assign PermutationsWithStreaming_mr_reset = reset;
  assign PermutationsWithStreaming_mr_io_in_0_Re = FFT_sr_v2_streaming_nrv_io_out_0_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_0_Im = FFT_sr_v2_streaming_nrv_io_out_0_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_1_Re = FFT_sr_v2_streaming_nrv_io_out_1_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_1_Im = FFT_sr_v2_streaming_nrv_io_out_1_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_2_Re = FFT_sr_v2_streaming_nrv_io_out_2_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_2_Im = FFT_sr_v2_streaming_nrv_io_out_2_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_3_Re = FFT_sr_v2_streaming_nrv_io_out_3_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_3_Im = FFT_sr_v2_streaming_nrv_io_out_3_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_4_Re = FFT_sr_v2_streaming_nrv_io_out_4_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_4_Im = FFT_sr_v2_streaming_nrv_io_out_4_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_5_Re = FFT_sr_v2_streaming_nrv_io_out_5_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_5_Im = FFT_sr_v2_streaming_nrv_io_out_5_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_6_Re = FFT_sr_v2_streaming_nrv_io_out_6_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_6_Im = FFT_sr_v2_streaming_nrv_io_out_6_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_7_Re = FFT_sr_v2_streaming_nrv_io_out_7_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_7_Im = FFT_sr_v2_streaming_nrv_io_out_7_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_en_0 = DFT_regdelays1_60; // @[FFTDesigns.scala 6489:37]
  assign PermutationsWithStreaming_mr_io_in_en_1 = Perm_regdelays1_1_0; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_2 = Perm_regdelays1_1_1; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_3 = Perm_regdelays1_1_2; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_4 = Perm_regdelays1_1_3; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_5 = Perm_regdelays1_1_4; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_6 = Perm_regdelays1_1_5; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_7 = Perm_regdelays1_1_6; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_8 = Perm_regdelays1_1_7; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_9 = Perm_regdelays1_1_8; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_10 = Perm_regdelays1_1_9; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_11 = Perm_regdelays1_1_10; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_12 = Perm_regdelays1_1_11; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_13 = Perm_regdelays1_1_12; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_14 = Perm_regdelays1_1_13; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_15 = Perm_regdelays1_1_14; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_16 = Perm_regdelays1_1_15; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_17 = Perm_regdelays1_1_16; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_18 = Perm_regdelays1_1_17; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_19 = Perm_regdelays1_1_18; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_20 = Perm_regdelays1_1_19; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_21 = Perm_regdelays1_1_20; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_22 = Perm_regdelays1_1_21; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_23 = Perm_regdelays1_1_22; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_24 = Perm_regdelays1_1_23; // @[FFTDesigns.scala 6513:51]
  assign PermutationsWithStreaming_mr_1_clock = clock;
  assign PermutationsWithStreaming_mr_1_reset = reset;
  assign PermutationsWithStreaming_mr_1_io_in_0_Re = DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_0_Im = DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_1_Re = DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_1_Im = DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_2_Re = DFT_r_v2_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_2_Im = DFT_r_v2_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_3_Re = DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_3_Im = DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_4_Re = DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_4_Im = DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_5_Re = DFT_r_v2_1_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_5_Im = DFT_r_v2_1_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_6_Re = DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_6_Im = DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_7_Re = DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_7_Im = DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_8_Re = DFT_r_v2_2_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_8_Im = DFT_r_v2_2_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_9_Re = DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_9_Im = DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_10_Re = DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_10_Im = DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_11_Re = DFT_r_v2_3_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_11_Im = DFT_r_v2_3_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_en_0 = DFT_regdelays2_3; // @[FFTDesigns.scala 6493:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_1 = Perm_regdelays1_2_0; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_2 = Perm_regdelays1_2_1; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_3 = Perm_regdelays1_2_2; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_4 = Perm_regdelays1_2_3; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_5 = Perm_regdelays1_2_4; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_6 = Perm_regdelays1_2_5; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_7 = Perm_regdelays1_2_6; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_8 = Perm_regdelays1_2_7; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_9 = Perm_regdelays1_2_8; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_10 = Perm_regdelays1_2_9; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_11 = Perm_regdelays1_2_10; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_12 = Perm_regdelays1_2_11; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_13 = Perm_regdelays1_2_12; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_14 = Perm_regdelays1_2_13; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_15 = Perm_regdelays1_2_14; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_16 = Perm_regdelays1_2_15; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_17 = Perm_regdelays1_2_16; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_18 = Perm_regdelays1_2_17; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_19 = Perm_regdelays1_2_18; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_20 = Perm_regdelays1_2_19; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_21 = Perm_regdelays1_2_20; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_22 = Perm_regdelays1_2_21; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_23 = Perm_regdelays1_2_22; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_24 = Perm_regdelays1_2_23; // @[FFTDesigns.scala 6515:51]
  assign TwiddleFactorsStreamed_mr_v2_clock = clock;
  assign TwiddleFactorsStreamed_mr_v2_reset = reset;
  assign TwiddleFactorsStreamed_mr_v2_io_in_0_Re = PermutationsWithStreaming_mr_io_out_0_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_0_Im = PermutationsWithStreaming_mr_io_out_0_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_1_Re = PermutationsWithStreaming_mr_io_out_1_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_1_Im = PermutationsWithStreaming_mr_io_out_1_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_2_Re = PermutationsWithStreaming_mr_io_out_2_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_2_Im = PermutationsWithStreaming_mr_io_out_2_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_3_Re = PermutationsWithStreaming_mr_io_out_3_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_3_Im = PermutationsWithStreaming_mr_io_out_3_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_4_Re = PermutationsWithStreaming_mr_io_out_4_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_4_Im = PermutationsWithStreaming_mr_io_out_4_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_5_Re = PermutationsWithStreaming_mr_io_out_5_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_5_Im = PermutationsWithStreaming_mr_io_out_5_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_6_Re = PermutationsWithStreaming_mr_io_out_6_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_6_Im = PermutationsWithStreaming_mr_io_out_6_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_7_Re = PermutationsWithStreaming_mr_io_out_7_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_7_Im = PermutationsWithStreaming_mr_io_out_7_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_8_Re = PermutationsWithStreaming_mr_io_out_8_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_8_Im = PermutationsWithStreaming_mr_io_out_8_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_9_Re = PermutationsWithStreaming_mr_io_out_9_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_9_Im = PermutationsWithStreaming_mr_io_out_9_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_10_Re = PermutationsWithStreaming_mr_io_out_10_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_10_Im = PermutationsWithStreaming_mr_io_out_10_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_11_Re = PermutationsWithStreaming_mr_io_out_11_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_11_Im = PermutationsWithStreaming_mr_io_out_11_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_en_0 = Perm_regdelays1_1_23; // @[FFTDesigns.scala 6524:33]
  assign TwiddleFactorsStreamed_mr_v2_io_in_en_1 = Twid_regdelays_0; // @[FFTDesigns.scala 6528:33]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_0 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_0 <= Perm_regdelays1_0_23; // @[FFTDesigns.scala 6534:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_1 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_1 <= DFT_regdelays1_0; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_2 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_2 <= DFT_regdelays1_1; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_3 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_3 <= DFT_regdelays1_2; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_4 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_4 <= DFT_regdelays1_3; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_5 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_5 <= DFT_regdelays1_4; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_6 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_6 <= DFT_regdelays1_5; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_7 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_7 <= DFT_regdelays1_6; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_8 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_8 <= DFT_regdelays1_7; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_9 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_9 <= DFT_regdelays1_8; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_10 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_10 <= DFT_regdelays1_9; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_11 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_11 <= DFT_regdelays1_10; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_12 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_12 <= DFT_regdelays1_11; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_13 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_13 <= DFT_regdelays1_12; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_14 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_14 <= DFT_regdelays1_13; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_15 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_15 <= DFT_regdelays1_14; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_16 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_16 <= DFT_regdelays1_15; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_17 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_17 <= DFT_regdelays1_16; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_18 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_18 <= DFT_regdelays1_17; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_19 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_19 <= DFT_regdelays1_18; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_20 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_20 <= DFT_regdelays1_19; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_21 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_21 <= DFT_regdelays1_20; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_22 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_22 <= DFT_regdelays1_21; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_23 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_23 <= DFT_regdelays1_22; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_24 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_24 <= DFT_regdelays1_23; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_25 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_25 <= DFT_regdelays1_24; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_26 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_26 <= DFT_regdelays1_25; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_27 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_27 <= DFT_regdelays1_26; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_28 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_28 <= DFT_regdelays1_27; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_29 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_29 <= DFT_regdelays1_28; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_30 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_30 <= DFT_regdelays1_29; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_31 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_31 <= DFT_regdelays1_30; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_32 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_32 <= DFT_regdelays1_31; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_33 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_33 <= DFT_regdelays1_32; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_34 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_34 <= DFT_regdelays1_33; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_35 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_35 <= DFT_regdelays1_34; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_36 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_36 <= DFT_regdelays1_35; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_37 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_37 <= DFT_regdelays1_36; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_38 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_38 <= DFT_regdelays1_37; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_39 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_39 <= DFT_regdelays1_38; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_40 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_40 <= DFT_regdelays1_39; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_41 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_41 <= DFT_regdelays1_40; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_42 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_42 <= DFT_regdelays1_41; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_43 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_43 <= DFT_regdelays1_42; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_44 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_44 <= DFT_regdelays1_43; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_45 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_45 <= DFT_regdelays1_44; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_46 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_46 <= DFT_regdelays1_45; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_47 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_47 <= DFT_regdelays1_46; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_48 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_48 <= DFT_regdelays1_47; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_49 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_49 <= DFT_regdelays1_48; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_50 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_50 <= DFT_regdelays1_49; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_51 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_51 <= DFT_regdelays1_50; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_52 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_52 <= DFT_regdelays1_51; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_53 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_53 <= DFT_regdelays1_52; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_54 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_54 <= DFT_regdelays1_53; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_55 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_55 <= DFT_regdelays1_54; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_56 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_56 <= DFT_regdelays1_55; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_57 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_57 <= DFT_regdelays1_56; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_58 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_58 <= DFT_regdelays1_57; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_59 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_59 <= DFT_regdelays1_58; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_60 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_60 <= DFT_regdelays1_59; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6475:35]
      DFT_regdelays2_0 <= 1'h0; // @[FFTDesigns.scala 6475:35]
    end else begin
      DFT_regdelays2_0 <= Twid_regdelays_1; // @[FFTDesigns.scala 6544:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6475:35]
      DFT_regdelays2_1 <= 1'h0; // @[FFTDesigns.scala 6475:35]
    end else begin
      DFT_regdelays2_1 <= DFT_regdelays2_0; // @[FFTDesigns.scala 6551:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6475:35]
      DFT_regdelays2_2 <= 1'h0; // @[FFTDesigns.scala 6475:35]
    end else begin
      DFT_regdelays2_2 <= DFT_regdelays2_1; // @[FFTDesigns.scala 6551:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6475:35]
      DFT_regdelays2_3 <= 1'h0; // @[FFTDesigns.scala 6475:35]
    end else begin
      DFT_regdelays2_3 <= DFT_regdelays2_2; // @[FFTDesigns.scala 6551:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6476:35]
      Twid_regdelays_0 <= 1'h0; // @[FFTDesigns.scala 6476:35]
    end else begin
      Twid_regdelays_0 <= Perm_regdelays1_1_23; // @[FFTDesigns.scala 6523:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6476:35]
      Twid_regdelays_1 <= 1'h0; // @[FFTDesigns.scala 6476:35]
    end else begin
      Twid_regdelays_1 <= Twid_regdelays_0; // @[FFTDesigns.scala 6527:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_0 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_0 <= io_in_ready; // @[FFTDesigns.scala 6484:37]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_1 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_1 <= Perm_regdelays1_0_0; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_2 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_2 <= Perm_regdelays1_0_1; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_3 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_3 <= Perm_regdelays1_0_2; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_4 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_4 <= Perm_regdelays1_0_3; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_5 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_5 <= Perm_regdelays1_0_4; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_6 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_6 <= Perm_regdelays1_0_5; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_7 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_7 <= Perm_regdelays1_0_6; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_8 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_8 <= Perm_regdelays1_0_7; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_9 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_9 <= Perm_regdelays1_0_8; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_10 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_10 <= Perm_regdelays1_0_9; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_11 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_11 <= Perm_regdelays1_0_10; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_12 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_12 <= Perm_regdelays1_0_11; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_13 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_13 <= Perm_regdelays1_0_12; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_14 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_14 <= Perm_regdelays1_0_13; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_15 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_15 <= Perm_regdelays1_0_14; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_16 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_16 <= Perm_regdelays1_0_15; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_17 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_17 <= Perm_regdelays1_0_16; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_18 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_18 <= Perm_regdelays1_0_17; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_19 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_19 <= Perm_regdelays1_0_18; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_20 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_20 <= Perm_regdelays1_0_19; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_21 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_21 <= Perm_regdelays1_0_20; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_22 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_22 <= Perm_regdelays1_0_21; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_23 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_23 <= Perm_regdelays1_0_22; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_0 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_0 <= DFT_regdelays1_60; // @[FFTDesigns.scala 6488:37]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_1 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_1 <= Perm_regdelays1_1_0; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_2 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_2 <= Perm_regdelays1_1_1; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_3 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_3 <= Perm_regdelays1_1_2; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_4 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_4 <= Perm_regdelays1_1_3; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_5 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_5 <= Perm_regdelays1_1_4; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_6 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_6 <= Perm_regdelays1_1_5; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_7 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_7 <= Perm_regdelays1_1_6; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_8 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_8 <= Perm_regdelays1_1_7; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_9 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_9 <= Perm_regdelays1_1_8; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_10 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_10 <= Perm_regdelays1_1_9; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_11 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_11 <= Perm_regdelays1_1_10; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_12 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_12 <= Perm_regdelays1_1_11; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_13 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_13 <= Perm_regdelays1_1_12; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_14 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_14 <= Perm_regdelays1_1_13; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_15 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_15 <= Perm_regdelays1_1_14; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_16 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_16 <= Perm_regdelays1_1_15; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_17 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_17 <= Perm_regdelays1_1_16; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_18 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_18 <= Perm_regdelays1_1_17; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_19 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_19 <= Perm_regdelays1_1_18; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_20 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_20 <= Perm_regdelays1_1_19; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_21 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_21 <= Perm_regdelays1_1_20; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_22 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_22 <= Perm_regdelays1_1_21; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_23 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_23 <= Perm_regdelays1_1_22; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_0 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_0 <= DFT_regdelays2_3; // @[FFTDesigns.scala 6492:37]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_1 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_1 <= Perm_regdelays1_2_0; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_2 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_2 <= Perm_regdelays1_2_1; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_3 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_3 <= Perm_regdelays1_2_2; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_4 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_4 <= Perm_regdelays1_2_3; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_5 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_5 <= Perm_regdelays1_2_4; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_6 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_6 <= Perm_regdelays1_2_5; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_7 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_7 <= Perm_regdelays1_2_6; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_8 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_8 <= Perm_regdelays1_2_7; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_9 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_9 <= Perm_regdelays1_2_8; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_10 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_10 <= Perm_regdelays1_2_9; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_11 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_11 <= Perm_regdelays1_2_10; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_12 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_12 <= Perm_regdelays1_2_11; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_13 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_13 <= Perm_regdelays1_2_12; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_14 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_14 <= Perm_regdelays1_2_13; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_15 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_15 <= Perm_regdelays1_2_14; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_16 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_16 <= Perm_regdelays1_2_15; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_17 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_17 <= Perm_regdelays1_2_16; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_18 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_18 <= Perm_regdelays1_2_17; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_19 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_19 <= Perm_regdelays1_2_18; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_20 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_20 <= Perm_regdelays1_2_19; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_21 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_21 <= Perm_regdelays1_2_20; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_22 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_22 <= Perm_regdelays1_2_21; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_23 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_23 <= Perm_regdelays1_2_22; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6478:33]
      out_regdelay <= 1'h0; // @[FFTDesigns.scala 6478:33]
    end else begin
      out_regdelay <= Perm_regdelays1_2_23; // @[FFTDesigns.scala 6554:20]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_0_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_0_Re <= PermutationsWithStreaming_mr_1_io_out_0_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_0_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_0_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_0_Im <= PermutationsWithStreaming_mr_1_io_out_0_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_0_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_1_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_1_Re <= PermutationsWithStreaming_mr_1_io_out_1_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_1_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_1_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_1_Im <= PermutationsWithStreaming_mr_1_io_out_1_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_1_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_2_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_2_Re <= PermutationsWithStreaming_mr_1_io_out_2_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_2_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_2_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_2_Im <= PermutationsWithStreaming_mr_1_io_out_2_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_2_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_3_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_3_Re <= PermutationsWithStreaming_mr_1_io_out_3_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_3_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_3_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_3_Im <= PermutationsWithStreaming_mr_1_io_out_3_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_3_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_4_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_4_Re <= PermutationsWithStreaming_mr_1_io_out_4_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_4_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_4_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_4_Im <= PermutationsWithStreaming_mr_1_io_out_4_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_4_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_5_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_5_Re <= PermutationsWithStreaming_mr_1_io_out_5_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_5_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_5_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_5_Im <= PermutationsWithStreaming_mr_1_io_out_5_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_5_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_6_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_6_Re <= PermutationsWithStreaming_mr_1_io_out_6_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_6_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_6_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_6_Im <= PermutationsWithStreaming_mr_1_io_out_6_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_6_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_7_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_7_Re <= PermutationsWithStreaming_mr_1_io_out_7_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_7_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_7_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_23) begin // @[FFTDesigns.scala 6555:49]
      results_7_Im <= PermutationsWithStreaming_mr_1_io_out_7_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_7_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DFT_regdelays1_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  DFT_regdelays1_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  DFT_regdelays1_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  DFT_regdelays1_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  DFT_regdelays1_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  DFT_regdelays1_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  DFT_regdelays1_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  DFT_regdelays1_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  DFT_regdelays1_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  DFT_regdelays1_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  DFT_regdelays1_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  DFT_regdelays1_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  DFT_regdelays1_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  DFT_regdelays1_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  DFT_regdelays1_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  DFT_regdelays1_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  DFT_regdelays1_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  DFT_regdelays1_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  DFT_regdelays1_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  DFT_regdelays1_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  DFT_regdelays1_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  DFT_regdelays1_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  DFT_regdelays1_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  DFT_regdelays1_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  DFT_regdelays1_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  DFT_regdelays1_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  DFT_regdelays1_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  DFT_regdelays1_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  DFT_regdelays1_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  DFT_regdelays1_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  DFT_regdelays1_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  DFT_regdelays1_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  DFT_regdelays1_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  DFT_regdelays1_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  DFT_regdelays1_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  DFT_regdelays1_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  DFT_regdelays1_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  DFT_regdelays1_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  DFT_regdelays1_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  DFT_regdelays1_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  DFT_regdelays1_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  DFT_regdelays1_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  DFT_regdelays1_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  DFT_regdelays1_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  DFT_regdelays1_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  DFT_regdelays1_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  DFT_regdelays1_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  DFT_regdelays1_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  DFT_regdelays1_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  DFT_regdelays1_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  DFT_regdelays1_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  DFT_regdelays1_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  DFT_regdelays1_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  DFT_regdelays1_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  DFT_regdelays1_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  DFT_regdelays1_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  DFT_regdelays1_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  DFT_regdelays1_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  DFT_regdelays1_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  DFT_regdelays1_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  DFT_regdelays1_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  DFT_regdelays2_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  DFT_regdelays2_1 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  DFT_regdelays2_2 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  DFT_regdelays2_3 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  Twid_regdelays_0 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  Twid_regdelays_1 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  Perm_regdelays1_0_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  Perm_regdelays1_0_1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  Perm_regdelays1_0_2 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  Perm_regdelays1_0_3 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  Perm_regdelays1_0_4 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  Perm_regdelays1_0_5 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  Perm_regdelays1_0_6 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  Perm_regdelays1_0_7 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  Perm_regdelays1_0_8 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  Perm_regdelays1_0_9 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  Perm_regdelays1_0_10 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  Perm_regdelays1_0_11 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  Perm_regdelays1_0_12 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  Perm_regdelays1_0_13 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  Perm_regdelays1_0_14 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  Perm_regdelays1_0_15 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  Perm_regdelays1_0_16 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  Perm_regdelays1_0_17 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  Perm_regdelays1_0_18 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  Perm_regdelays1_0_19 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  Perm_regdelays1_0_20 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  Perm_regdelays1_0_21 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  Perm_regdelays1_0_22 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  Perm_regdelays1_0_23 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  Perm_regdelays1_1_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  Perm_regdelays1_1_1 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  Perm_regdelays1_1_2 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  Perm_regdelays1_1_3 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  Perm_regdelays1_1_4 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  Perm_regdelays1_1_5 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  Perm_regdelays1_1_6 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  Perm_regdelays1_1_7 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  Perm_regdelays1_1_8 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  Perm_regdelays1_1_9 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  Perm_regdelays1_1_10 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  Perm_regdelays1_1_11 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  Perm_regdelays1_1_12 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  Perm_regdelays1_1_13 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  Perm_regdelays1_1_14 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  Perm_regdelays1_1_15 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  Perm_regdelays1_1_16 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  Perm_regdelays1_1_17 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  Perm_regdelays1_1_18 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  Perm_regdelays1_1_19 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  Perm_regdelays1_1_20 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  Perm_regdelays1_1_21 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  Perm_regdelays1_1_22 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  Perm_regdelays1_1_23 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  Perm_regdelays1_2_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  Perm_regdelays1_2_1 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  Perm_regdelays1_2_2 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  Perm_regdelays1_2_3 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  Perm_regdelays1_2_4 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  Perm_regdelays1_2_5 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  Perm_regdelays1_2_6 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  Perm_regdelays1_2_7 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  Perm_regdelays1_2_8 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  Perm_regdelays1_2_9 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  Perm_regdelays1_2_10 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  Perm_regdelays1_2_11 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  Perm_regdelays1_2_12 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  Perm_regdelays1_2_13 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  Perm_regdelays1_2_14 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  Perm_regdelays1_2_15 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  Perm_regdelays1_2_16 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  Perm_regdelays1_2_17 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  Perm_regdelays1_2_18 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  Perm_regdelays1_2_19 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  Perm_regdelays1_2_20 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  Perm_regdelays1_2_21 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  Perm_regdelays1_2_22 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  Perm_regdelays1_2_23 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  out_regdelay = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  results_0_Re = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  results_0_Im = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  results_1_Re = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  results_1_Im = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  results_2_Re = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  results_2_Im = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  results_3_Re = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  results_3_Im = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  results_4_Re = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  results_4_Im = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  results_5_Re = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  results_5_Im = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  results_6_Re = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  results_6_Im = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  results_7_Re = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  results_7_Im = _RAND_155[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

