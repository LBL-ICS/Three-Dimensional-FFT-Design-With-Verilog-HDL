module full_subber(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[Arithmetic.scala 72:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[Arithmetic.scala 72:34]
  wire [8:0] result = _result_T_2[8:0]; // @[Arithmetic.scala 71:22 72:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 73:23]
  assign io_out_c = result[8]; // @[Arithmetic.scala 74:23]
endmodule
module twoscomplement(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _x_T = ~io_in; // @[Arithmetic.scala 28:16]
  assign io_out = 8'h1 + _x_T; // @[Arithmetic.scala 28:14]
endmodule
module full_adder(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 58:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 58:34]
  wire [24:0] result = _result_T_1[24:0]; // @[Arithmetic.scala 57:22 58:12]
  assign io_out_s = result[23:0]; // @[Arithmetic.scala 59:23]
  assign io_out_c = result[24]; // @[Arithmetic.scala 60:23]
endmodule
module twoscomplement_1(
  input  [23:0] io_in,
  output [23:0] io_out
);
  wire [23:0] _x_T = ~io_in; // @[Arithmetic.scala 28:16]
  assign io_out = 24'h1 + _x_T; // @[Arithmetic.scala 28:14]
endmodule
module shifter(
  input  [23:0] io_in_a,
  input  [4:0]  io_in_b,
  output [23:0] io_out_s
);
  wire [23:0] _result_T = io_in_a >> io_in_b; // @[Arithmetic.scala 42:25]
  wire [54:0] _GEN_0 = {{31'd0}, _result_T}; // @[Arithmetic.scala 41:26 42:14 44:14]
  assign io_out_s = _GEN_0[23:0]; // @[Arithmetic.scala 39:22]
endmodule
module leadingOneDetector(
  input  [23:0] io_in,
  output [4:0]  io_out
);
  wire [1:0] _hotValue_T = io_in[1] ? 2'h2 : 2'h1; // @[Mux.scala 47:70]
  wire [1:0] _hotValue_T_1 = io_in[2] ? 2'h3 : _hotValue_T; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_2 = io_in[3] ? 3'h4 : {{1'd0}, _hotValue_T_1}; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_3 = io_in[4] ? 3'h5 : _hotValue_T_2; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_4 = io_in[5] ? 3'h6 : _hotValue_T_3; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_5 = io_in[6] ? 3'h7 : _hotValue_T_4; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_6 = io_in[7] ? 4'h8 : {{1'd0}, _hotValue_T_5}; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_7 = io_in[8] ? 4'h9 : _hotValue_T_6; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_8 = io_in[9] ? 4'ha : _hotValue_T_7; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_9 = io_in[10] ? 4'hb : _hotValue_T_8; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_10 = io_in[11] ? 4'hc : _hotValue_T_9; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_11 = io_in[12] ? 4'hd : _hotValue_T_10; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_12 = io_in[13] ? 4'he : _hotValue_T_11; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_13 = io_in[14] ? 4'hf : _hotValue_T_12; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_14 = io_in[15] ? 5'h10 : {{1'd0}, _hotValue_T_13}; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_15 = io_in[16] ? 5'h11 : _hotValue_T_14; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_16 = io_in[17] ? 5'h12 : _hotValue_T_15; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_17 = io_in[18] ? 5'h13 : _hotValue_T_16; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_18 = io_in[19] ? 5'h14 : _hotValue_T_17; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_19 = io_in[20] ? 5'h15 : _hotValue_T_18; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_20 = io_in[21] ? 5'h16 : _hotValue_T_19; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_21 = io_in[22] ? 5'h17 : _hotValue_T_20; // @[Mux.scala 47:70]
  assign io_out = io_in[23] ? 5'h18 : _hotValue_T_21; // @[Mux.scala 47:70]
endmodule
module FP_adder(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 76:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 76:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 76:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 76:24]
  wire [7:0] complement_io_in; // @[FPArithmetic.scala 82:28]
  wire [7:0] complement_io_out; // @[FPArithmetic.scala 82:28]
  wire [23:0] adder_io_in_a; // @[FPArithmetic.scala 86:23]
  wire [23:0] adder_io_in_b; // @[FPArithmetic.scala 86:23]
  wire [23:0] adder_io_out_s; // @[FPArithmetic.scala 86:23]
  wire  adder_io_out_c; // @[FPArithmetic.scala 86:23]
  wire [23:0] complementN_0_io_in; // @[FPArithmetic.scala 92:31]
  wire [23:0] complementN_0_io_out; // @[FPArithmetic.scala 92:31]
  wire [23:0] complementN_1_io_in; // @[FPArithmetic.scala 94:31]
  wire [23:0] complementN_1_io_out; // @[FPArithmetic.scala 94:31]
  wire [23:0] shifter_io_in_a; // @[FPArithmetic.scala 98:25]
  wire [4:0] shifter_io_in_b; // @[FPArithmetic.scala 98:25]
  wire [23:0] shifter_io_out_s; // @[FPArithmetic.scala 98:25]
  wire [23:0] complementN_2_io_in; // @[FPArithmetic.scala 143:31]
  wire [23:0] complementN_2_io_out; // @[FPArithmetic.scala 143:31]
  wire [23:0] leadingOneFinder_io_in; // @[FPArithmetic.scala 163:34]
  wire [4:0] leadingOneFinder_io_out; // @[FPArithmetic.scala 163:34]
  wire [7:0] subber2_io_in_a; // @[FPArithmetic.scala 165:25]
  wire [7:0] subber2_io_in_b; // @[FPArithmetic.scala 165:25]
  wire [7:0] subber2_io_out_s; // @[FPArithmetic.scala 165:25]
  wire  subber2_io_out_c; // @[FPArithmetic.scala 165:25]
  wire  sign_0 = io_in_a[31]; // @[FPArithmetic.scala 38:23]
  wire  sign_1 = io_in_b[31]; // @[FPArithmetic.scala 39:23]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 43:62]
  wire [8:0] _GEN_31 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 43:34]
  wire [8:0] _GEN_0 = _GEN_31 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 43:68 44:14 46:14]
  wire [8:0] _GEN_32 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 48:34]
  wire [8:0] _GEN_1 = _GEN_32 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 48:68 49:14 51:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 56:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 57:23]
  wire [23:0] whole_frac_0 = {1'h1,frac_0}; // @[FPArithmetic.scala 61:26]
  wire [23:0] whole_frac_1 = {1'h1,frac_1}; // @[FPArithmetic.scala 62:26]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 42:19]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 42:19]
  wire [7:0] out_exp = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 104:34 105:15 115:15]
  wire [7:0] sub_exp = subber_io_out_c ? complement_io_out : subber_io_out_s; // @[FPArithmetic.scala 104:34 106:15 116:15]
  wire  out_s = subber_io_out_c ? sign_1 : sign_0; // @[FPArithmetic.scala 104:34 107:13 117:13]
  wire [22:0] out_frac = subber_io_out_c ? frac_1 : frac_0; // @[FPArithmetic.scala 104:34 108:16 118:16]
  wire [23:0] _GEN_8 = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 104:34 112:21 87:19]
  wire [23:0] _GEN_9 = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 104:34 88:19 122:21]
  wire  _new_s_T = ~adder_io_out_c; // @[FPArithmetic.scala 138:15]
  wire  _D_T_1 = sign_0 ^ sign_1; // @[FPArithmetic.scala 151:39]
  wire  D = _new_s_T | sign_0 ^ sign_1; // @[FPArithmetic.scala 151:28]
  wire  E = _new_s_T & ~adder_io_out_s[23] | _new_s_T & ~_D_T_1 | adder_io_out_c & adder_io_out_s[23] & _D_T_1; // @[FPArithmetic.scala 154:99]
  wire  _GEN_25 = sub_exp >= 8'h17 ? out_s : ~adder_io_out_c & sign_0 | sign_0 & sign_1 | ~adder_io_out_c & sign_1; // @[FPArithmetic.scala 138:11 173:39 174:13]
  wire  new_s = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 1'h0 : _GEN_25; // @[FPArithmetic.scala 169:62 170:13]
  wire [23:0] adder_result = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 157:18 158:47 159:20]
  wire [4:0] _subber2_io_in_b_T_1 = 5'h18 - leadingOneFinder_io_out; // @[FPArithmetic.scala 167:42]
  wire [8:0] _GEN_33 = {{1'd0}, out_exp}; // @[FPArithmetic.scala 181:20]
  wire [23:0] _new_out_frac_T_2 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 183:51]
  wire [7:0] _new_out_exp_T_3 = out_exp + 8'h1; // @[FPArithmetic.scala 185:32]
  wire [8:0] _GEN_13 = _GEN_33 == _T_2 ? _T_2 : {{1'd0}, _new_out_exp_T_3}; // @[FPArithmetic.scala 181:56 182:21 185:21]
  wire [23:0] _GEN_14 = _GEN_33 == _T_2 ? _new_out_frac_T_2 : {{1'd0}, adder_result[23:1]}; // @[FPArithmetic.scala 181:56 183:22 186:22]
  wire [53:0] _GEN_2 = {{31'd0}, adder_result[22:0]}; // @[FPArithmetic.scala 197:57]
  wire [53:0] _new_out_frac_T_7 = _GEN_2 << _subber2_io_in_b_T_1; // @[FPArithmetic.scala 197:57]
  wire [7:0] _GEN_15 = subber2_io_out_c ? 8'h1 : subber2_io_out_s; // @[FPArithmetic.scala 192:39 193:23 196:23]
  wire [53:0] _GEN_16 = subber2_io_out_c ? 54'h400000 : _new_out_frac_T_7; // @[FPArithmetic.scala 192:39 194:24 197:24]
  wire [7:0] _GEN_17 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:0
    ]) ? 8'h0 : _GEN_15; // @[FPArithmetic.scala 189:141 190:21]
  wire [53:0] _GEN_18 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:
    0]) ? 54'h0 : _GEN_16; // @[FPArithmetic.scala 189:141 139:18]
  wire [7:0] _GEN_19 = D ? _GEN_17 : 8'h0; // @[FPArithmetic.scala 140:17 188:26]
  wire [53:0] _GEN_20 = D ? _GEN_18 : 54'h0; // @[FPArithmetic.scala 139:18 188:26]
  wire [8:0] _GEN_21 = ~D ? _GEN_13 : {{1'd0}, _GEN_19}; // @[FPArithmetic.scala 180:26]
  wire [53:0] _GEN_22 = ~D ? {{30'd0}, _GEN_14} : _GEN_20; // @[FPArithmetic.scala 180:26]
  wire [8:0] _GEN_23 = E ? {{1'd0}, out_exp} : _GEN_21; // @[FPArithmetic.scala 177:26 178:19]
  wire [53:0] _GEN_24 = E ? {{31'd0}, adder_result[22:0]} : _GEN_22; // @[FPArithmetic.scala 177:26 179:20]
  wire [53:0] _GEN_26 = sub_exp >= 8'h17 ? {{31'd0}, out_frac} : _GEN_24; // @[FPArithmetic.scala 173:39 175:20]
  wire [8:0] _GEN_27 = sub_exp >= 8'h17 ? {{1'd0}, out_exp} : _GEN_23; // @[FPArithmetic.scala 173:39 176:19]
  wire [8:0] _GEN_29 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 9'h0 : _GEN_27; // @[FPArithmetic.scala 169:62 171:19]
  wire [53:0] _GEN_30 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 54'h0 : _GEN_26; // @[FPArithmetic.scala 169:62 172:20]
  reg [31:0] reg_out_s; // @[FPArithmetic.scala 201:28]
  wire [7:0] new_out_exp = _GEN_29[7:0]; // @[FPArithmetic.scala 137:27]
  wire [22:0] new_out_frac = _GEN_30[22:0]; // @[FPArithmetic.scala 136:28]
  wire [31:0] _reg_out_s_T_1 = {new_s,new_out_exp,new_out_frac}; // @[FPArithmetic.scala 203:39]
  full_subber subber ( // @[FPArithmetic.scala 76:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complement ( // @[FPArithmetic.scala 82:28]
    .io_in(complement_io_in),
    .io_out(complement_io_out)
  );
  full_adder adder ( // @[FPArithmetic.scala 86:23]
    .io_in_a(adder_io_in_a),
    .io_in_b(adder_io_in_b),
    .io_out_s(adder_io_out_s),
    .io_out_c(adder_io_out_c)
  );
  twoscomplement_1 complementN_0 ( // @[FPArithmetic.scala 92:31]
    .io_in(complementN_0_io_in),
    .io_out(complementN_0_io_out)
  );
  twoscomplement_1 complementN_1 ( // @[FPArithmetic.scala 94:31]
    .io_in(complementN_1_io_in),
    .io_out(complementN_1_io_out)
  );
  shifter shifter ( // @[FPArithmetic.scala 98:25]
    .io_in_a(shifter_io_in_a),
    .io_in_b(shifter_io_in_b),
    .io_out_s(shifter_io_out_s)
  );
  twoscomplement_1 complementN_2 ( // @[FPArithmetic.scala 143:31]
    .io_in(complementN_2_io_in),
    .io_out(complementN_2_io_out)
  );
  leadingOneDetector leadingOneFinder ( // @[FPArithmetic.scala 163:34]
    .io_in(leadingOneFinder_io_in),
    .io_out(leadingOneFinder_io_out)
  );
  full_subber subber2 ( // @[FPArithmetic.scala 165:25]
    .io_in_a(subber2_io_in_a),
    .io_in_b(subber2_io_in_b),
    .io_out_s(subber2_io_out_s),
    .io_out_c(subber2_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FPArithmetic.scala 205:14]
  assign subber_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 42:19]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 42:19]
  assign complement_io_in = subber_io_out_s; // @[FPArithmetic.scala 83:22]
  assign adder_io_in_a = sign_0 & ~sign_1 ? complementN_0_io_out : _GEN_8; // @[FPArithmetic.scala 127:45 128:21]
  assign adder_io_in_b = sign_1 & ~sign_0 ? complementN_1_io_out : _GEN_9; // @[FPArithmetic.scala 131:45 132:21]
  assign complementN_0_io_in = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 104:34 112:21 87:19]
  assign complementN_1_io_in = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 104:34 88:19 122:21]
  assign shifter_io_in_a = subber_io_out_c ? whole_frac_0 : whole_frac_1; // @[FPArithmetic.scala 104:34 109:23 119:23]
  assign shifter_io_in_b = sub_exp[4:0];
  assign complementN_2_io_in = adder_io_out_s; // @[FPArithmetic.scala 144:25]
  assign leadingOneFinder_io_in = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 157:18 158:47 159:20]
  assign subber2_io_in_a = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 104:34 105:15 115:15]
  assign subber2_io_in_b = {{3'd0}, _subber2_io_in_b_T_1}; // @[FPArithmetic.scala 167:21]
  always @(posedge clock) begin
    if (reset) begin // @[FPArithmetic.scala 201:28]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 201:28]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FPArithmetic.scala 203:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_out_s = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexAdder(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_adder_clock; // @[FPComplex.scala 21:25]
  wire  FP_adder_reset; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 21:25]
  wire  FP_adder_1_clock; // @[FPComplex.scala 21:25]
  wire  FP_adder_1_reset; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_in_a; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_in_b; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_out_s; // @[FPComplex.scala 21:25]
  FP_adder FP_adder ( // @[FPComplex.scala 21:25]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_adder FP_adder_1 ( // @[FPComplex.scala 21:25]
    .clock(FP_adder_1_clock),
    .reset(FP_adder_1_reset),
    .io_in_a(FP_adder_1_io_in_a),
    .io_in_b(FP_adder_1_io_in_b),
    .io_out_s(FP_adder_1_io_out_s)
  );
  assign io_out_s_Re = FP_adder_io_out_s; // @[FPComplex.scala 28:17]
  assign io_out_s_Im = FP_adder_1_io_out_s; // @[FPComplex.scala 29:17]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = io_in_a_Re; // @[FPComplex.scala 24:23]
  assign FP_adder_io_in_b = io_in_b_Re; // @[FPComplex.scala 25:23]
  assign FP_adder_1_clock = clock;
  assign FP_adder_1_reset = reset;
  assign FP_adder_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 26:23]
  assign FP_adder_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 27:23]
endmodule
module FP_subber(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_clock; // @[FPArithmetic.scala 414:26]
  wire  FP_adder_reset; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_in_a; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_in_b; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_out_s; // @[FPArithmetic.scala 414:26]
  wire  _adjusted_in_b_T_1 = ~io_in_b[31]; // @[FPArithmetic.scala 417:23]
  FP_adder FP_adder ( // @[FPArithmetic.scala 414:26]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  assign io_out_s = FP_adder_io_out_s; // @[FPArithmetic.scala 420:14]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = io_in_a; // @[FPArithmetic.scala 418:22]
  assign FP_adder_io_in_b = {_adjusted_in_b_T_1,io_in_b[30:0]}; // @[FPArithmetic.scala 417:39]
endmodule
module FPComplexSub(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_subber_clock; // @[FPComplex.scala 78:25]
  wire  FP_subber_reset; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 78:25]
  wire  FP_subber_1_clock; // @[FPComplex.scala 78:25]
  wire  FP_subber_1_reset; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_in_a; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_in_b; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_out_s; // @[FPComplex.scala 78:25]
  FP_subber FP_subber ( // @[FPComplex.scala 78:25]
    .clock(FP_subber_clock),
    .reset(FP_subber_reset),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_subber FP_subber_1 ( // @[FPComplex.scala 78:25]
    .clock(FP_subber_1_clock),
    .reset(FP_subber_1_reset),
    .io_in_a(FP_subber_1_io_in_a),
    .io_in_b(FP_subber_1_io_in_b),
    .io_out_s(FP_subber_1_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 85:17]
  assign io_out_s_Im = FP_subber_1_io_out_s; // @[FPComplex.scala 86:17]
  assign FP_subber_clock = clock;
  assign FP_subber_reset = reset;
  assign FP_subber_io_in_a = io_in_a_Re; // @[FPComplex.scala 81:24]
  assign FP_subber_io_in_b = io_in_b_Re; // @[FPComplex.scala 82:24]
  assign FP_subber_1_clock = clock;
  assign FP_subber_1_reset = reset;
  assign FP_subber_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 83:24]
  assign FP_subber_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 84:24]
endmodule
module FPComplexMultiAdder(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  assign io_out_Re = io_in_0_Re; // @[FPComplex.scala 474:14]
  assign io_out_Im = io_in_0_Im; // @[FPComplex.scala 474:14]
endmodule
module cmplx_adj(
  input  [31:0] io_in_Re,
  input  [31:0] io_in_Im,
  input  [7:0]  io_in_adj,
  input         io_is_neg,
  input         io_is_flip,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  wire  sign_0 = io_in_Re[31]; // @[FFTDesigns.scala 3510:24]
  wire  sign_1 = io_in_Im[31]; // @[FFTDesigns.scala 3511:24]
  wire [7:0] exp_0 = io_in_Re[30:23]; // @[FFTDesigns.scala 3513:23]
  wire [7:0] exp_1 = io_in_Im[30:23]; // @[FFTDesigns.scala 3514:23]
  wire [22:0] frac_0 = io_in_Re[22:0]; // @[FFTDesigns.scala 3516:24]
  wire [22:0] frac_1 = io_in_Im[22:0]; // @[FFTDesigns.scala 3517:24]
  wire  new_sign_0 = io_is_neg ? ~sign_0 : sign_0; // @[FFTDesigns.scala 3519:20 3520:19 3523:19]
  wire  new_sign_1 = io_is_neg ? ~sign_1 : sign_1; // @[FFTDesigns.scala 3519:20 3521:19 3524:19]
  wire [7:0] _new_exp_0_T_1 = exp_0 - io_in_adj; // @[FFTDesigns.scala 3528:28]
  wire [7:0] new_exp_0 = exp_0 != 8'h0 ? _new_exp_0_T_1 : exp_0; // @[FFTDesigns.scala 3527:25 3528:18 3530:18]
  wire [7:0] _new_exp_1_T_1 = exp_1 - io_in_adj; // @[FFTDesigns.scala 3533:28]
  wire [7:0] new_exp_1 = exp_1 != 8'h0 ? _new_exp_1_T_1 : exp_1; // @[FFTDesigns.scala 3532:26 3533:18 3535:18]
  wire  _io_out_Re_T = ~new_sign_1; // @[FFTDesigns.scala 3539:21]
  wire [31:0] _io_out_Re_T_2 = {_io_out_Re_T,new_exp_1,frac_1}; // @[FFTDesigns.scala 3539:49]
  wire [31:0] _io_out_Im_T_1 = {new_sign_0,new_exp_0,frac_0}; // @[FFTDesigns.scala 3540:48]
  wire [31:0] _io_out_Im_T_3 = {new_sign_1,new_exp_1,frac_1}; // @[FFTDesigns.scala 3543:48]
  assign io_out_Re = io_is_flip ? _io_out_Re_T_2 : _io_out_Im_T_1; // @[FFTDesigns.scala 3538:21 3539:17 3542:17]
  assign io_out_Im = io_is_flip ? _io_out_Im_T_1 : _io_out_Im_T_3; // @[FFTDesigns.scala 3538:21 3540:17 3543:17]
endmodule
module FPComplexMult_reducable_v2(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 333:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 333:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 333:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 333:33]
  reg [31:0] result_0_Re; // @[FPComplex.scala 344:31]
  reg [31:0] result_0_Im; // @[FPComplex.scala 344:31]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 333:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  assign io_out_s_Re = result_0_Re; // @[FPComplex.scala 353:20]
  assign io_out_s_Im = result_0_Im; // @[FPComplex.scala 353:20]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 334:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 334:24]
  assign cmplx_adj_io_in_adj = 8'h1; // @[FPComplex.scala 337:30]
  assign cmplx_adj_io_is_neg = 1'h1; // @[FPComplex.scala 339:32]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FPComplex.scala 335:29]
  always @(posedge clock) begin
    if (reset) begin // @[FPComplex.scala 344:31]
      result_0_Re <= 32'h0; // @[FPComplex.scala 344:31]
    end else begin
      result_0_Re <= cmplx_adj_io_out_Re; // @[FPComplex.scala 347:25]
    end
    if (reset) begin // @[FPComplex.scala 344:31]
      result_0_Im <= 32'h0; // @[FPComplex.scala 344:31]
    end else begin
      result_0_Im <= cmplx_adj_io_out_Im; // @[FPComplex.scala 347:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  result_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  result_0_Im = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multiplier(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[Arithmetic.scala 84:23]
endmodule
module full_adder_4(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 58:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 58:34]
  wire [8:0] result = _result_T_1[8:0]; // @[Arithmetic.scala 57:22 58:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 59:23]
endmodule
module FP_multiplier(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] multiplier_io_in_a; // @[FPArithmetic.scala 488:28]
  wire [23:0] multiplier_io_in_b; // @[FPArithmetic.scala 488:28]
  wire [47:0] multiplier_io_out_s; // @[FPArithmetic.scala 488:28]
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 493:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 493:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 493:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 493:24]
  wire [7:0] complementN_io_in; // @[FPArithmetic.scala 499:29]
  wire [7:0] complementN_io_out; // @[FPArithmetic.scala 499:29]
  wire [7:0] adderN_io_in_a; // @[FPArithmetic.scala 503:24]
  wire [7:0] adderN_io_in_b; // @[FPArithmetic.scala 503:24]
  wire [7:0] adderN_io_out_s; // @[FPArithmetic.scala 503:24]
  wire  s_0 = io_in_a[31]; // @[FPArithmetic.scala 453:20]
  wire  s_1 = io_in_b[31]; // @[FPArithmetic.scala 454:20]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 458:62]
  wire [8:0] _GEN_13 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 458:34]
  wire [8:0] _GEN_0 = _GEN_13 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 458:68 459:14 461:14]
  wire [8:0] _GEN_14 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 463:34]
  wire [8:0] _GEN_1 = _GEN_14 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 463:68 464:14 466:14]
  wire [22:0] exp_check_0 = {{15'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 469:25 470:18]
  wire [22:0] _cond_holder_T_1 = exp_check_0 + 23'h1; // @[FPArithmetic.scala 474:34]
  wire [22:0] exp_check_1 = {{15'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 469:25 471:18]
  wire [22:0] _cond_holder_T_3 = 23'h7f - exp_check_1; // @[FPArithmetic.scala 474:80]
  wire [22:0] _cond_holder_T_4 = ~_cond_holder_T_3; // @[FPArithmetic.scala 474:42]
  wire [22:0] _cond_holder_T_6 = _cond_holder_T_1 + _cond_holder_T_4; // @[FPArithmetic.scala 474:40]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 478:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 479:23]
  wire  new_s = s_0 ^ s_1; // @[FPArithmetic.scala 510:19]
  wire [7:0] _new_exp_T_1 = adderN_io_out_s + 8'h1; // @[FPArithmetic.scala 521:34]
  wire [22:0] _cond_holder_T_8 = exp_check_0 + 23'h2; // @[FPArithmetic.scala 523:36]
  wire [22:0] _cond_holder_T_13 = _cond_holder_T_8 + _cond_holder_T_4; // @[FPArithmetic.scala 523:42]
  wire [23:0] _new_mant_T_2 = {multiplier_io_out_s[46:24], 1'h0}; // @[FPArithmetic.scala 529:73]
  wire [7:0] _GEN_2 = multiplier_io_out_s[47] ? _new_exp_T_1 : adderN_io_out_s; // @[FPArithmetic.scala 520:60 521:15 526:15]
  wire [22:0] cond_holder = multiplier_io_out_s[47] ? _cond_holder_T_13 : _cond_holder_T_6; // @[FPArithmetic.scala 520:60 523:19 528:19]
  wire [23:0] _GEN_5 = multiplier_io_out_s[47] ? {{1'd0}, multiplier_io_out_s[46:24]} : _new_mant_T_2; // @[FPArithmetic.scala 520:60 524:16 529:16]
  reg [31:0] reg_out_s; // @[FPArithmetic.scala 531:28]
  wire [22:0] _T_12 = ~cond_holder; // @[FPArithmetic.scala 533:51]
  wire [22:0] _T_14 = 23'h1 + _T_12; // @[FPArithmetic.scala 533:49]
  wire [22:0] _GEN_15 = {{14'd0}, _T_2}; // @[FPArithmetic.scala 533:42]
  wire [8:0] _GEN_6 = cond_holder > _GEN_15 ? _T_2 : {{1'd0}, _GEN_2}; // @[FPArithmetic.scala 538:61 539:15]
  wire [8:0] _GEN_9 = _GEN_15 >= _T_14 ? 9'h1 : _GEN_6; // @[FPArithmetic.scala 533:67 534:15]
  wire [7:0] new_exp = _GEN_9[7:0]; // @[FPArithmetic.scala 513:23]
  wire [23:0] _new_mant_T_4 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 540:45]
  wire [23:0] _GEN_7 = cond_holder > _GEN_15 ? _new_mant_T_4 : _GEN_5; // @[FPArithmetic.scala 538:61 540:16]
  wire [23:0] _GEN_10 = _GEN_15 >= _T_14 ? 24'h400000 : _GEN_7; // @[FPArithmetic.scala 533:67 535:16]
  wire [22:0] new_mant = _GEN_10[22:0]; // @[FPArithmetic.scala 515:24]
  wire [31:0] _reg_out_s_T_1 = {new_s,new_exp,new_mant}; // @[FPArithmetic.scala 536:37]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 457:19]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 457:19]
  multiplier multiplier ( // @[FPArithmetic.scala 488:28]
    .io_in_a(multiplier_io_in_a),
    .io_in_b(multiplier_io_in_b),
    .io_out_s(multiplier_io_out_s)
  );
  full_subber subber ( // @[FPArithmetic.scala 493:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complementN ( // @[FPArithmetic.scala 499:29]
    .io_in(complementN_io_in),
    .io_out(complementN_io_out)
  );
  full_adder_4 adderN ( // @[FPArithmetic.scala 503:24]
    .io_in_a(adderN_io_in_a),
    .io_in_b(adderN_io_in_b),
    .io_out_s(adderN_io_out_s)
  );
  assign io_out_s = reg_out_s; // @[FPArithmetic.scala 548:14]
  assign multiplier_io_in_a = {1'h1,frac_0}; // @[FPArithmetic.scala 483:24]
  assign multiplier_io_in_b = {1'h1,frac_1}; // @[FPArithmetic.scala 484:24]
  assign subber_io_in_a = 8'h7f; // @[FPArithmetic.scala 494:20]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 457:19]
  assign complementN_io_in = subber_io_out_s; // @[FPArithmetic.scala 500:23]
  assign adderN_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 457:19]
  assign adderN_io_in_b = complementN_io_out; // @[FPArithmetic.scala 505:20]
  always @(posedge clock) begin
    if (reset) begin // @[FPArithmetic.scala 531:28]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 531:28]
    end else if (exp_0 == 8'h0 | exp_1 == 8'h0) begin // @[FPArithmetic.scala 543:43]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 544:17]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FPArithmetic.scala 546:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_out_s = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMult_reducable_v2_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 293:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 293:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 293:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 293:33]
  wire  FP_multiplier_clock; // @[FPComplex.scala 321:29]
  wire  FP_multiplier_reset; // @[FPComplex.scala 321:29]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 321:29]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 321:29]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 321:29]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 321:29]
  wire  FP_multiplier_1_reset; // @[FPComplex.scala 321:29]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 321:29]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 321:29]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 321:29]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 293:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 321:29]
    .clock(FP_multiplier_clock),
    .reset(FP_multiplier_reset),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 321:29]
    .clock(FP_multiplier_1_clock),
    .reset(FP_multiplier_1_reset),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  assign io_out_s_Re = FP_multiplier_io_out_s; // @[FPComplex.scala 328:21]
  assign io_out_s_Im = FP_multiplier_1_io_out_s; // @[FPComplex.scala 329:21]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 294:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 294:24]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FPComplex.scala 318:30]
  assign cmplx_adj_io_is_neg = 1'h0; // @[FPComplex.scala 319:30]
  assign cmplx_adj_io_is_flip = 1'h1; // @[FPComplex.scala 295:29]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_reset = reset;
  assign FP_multiplier_io_in_a = cmplx_adj_io_out_Re; // @[FPComplex.scala 324:29]
  assign FP_multiplier_io_in_b = 32'hbf5db3d6; // @[FPComplex.scala 325:29]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_reset = reset;
  assign FP_multiplier_1_io_in_a = cmplx_adj_io_out_Im; // @[FPComplex.scala 326:29]
  assign FP_multiplier_1_io_in_b = 32'hbf5db3d6; // @[FPComplex.scala 327:29]
endmodule
module DFT_r_v2(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  FPComplexAdder_clock; // @[FFTDesigns.scala 258:34]
  wire  FPComplexAdder_reset; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_a_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_a_Im; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_b_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_b_Im; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 258:34]
  wire  FPComplexSub_clock; // @[FFTDesigns.scala 261:34]
  wire  FPComplexSub_reset; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_a_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_a_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_b_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_b_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_out_s_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_out_s_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexMultiAdder_io_in_0_Re; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_in_0_Im; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 275:36]
  wire  FPComplexMult_reducable_v2_clock; // @[FFTDesigns.scala 294:39]
  wire  FPComplexMult_reducable_v2_reset; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Re; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Im; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 294:39]
  wire  FPComplexMult_reducable_v2_1_clock; // @[FFTDesigns.scala 297:39]
  wire  FPComplexMult_reducable_v2_1_reset; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Re; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Im; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 297:39]
  wire  FPComplexAdder_reducable_clock; // @[FFTDesigns.scala 338:34]
  wire  FPComplexAdder_reducable_reset; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_a_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_a_Im; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_b_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_b_Im; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_out_s_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_out_s_Im; // @[FFTDesigns.scala 338:34]
  wire  FPComplexSub_reducable_clock; // @[FFTDesigns.scala 341:34]
  wire  FPComplexSub_reducable_reset; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_a_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_a_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_b_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_b_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_out_s_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_out_s_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_in_0_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_in_0_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_out_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_out_Im; // @[FFTDesigns.scala 394:29]
  wire  FPComplexAdder_1_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_1_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_2_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_2_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_3_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_3_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  reg [31:0] initial_layer_out_0_0_Re; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_0_0_Im; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_1_0_Re; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_1_0_Im; // @[FFTDesigns.scala 276:84]
  reg [31:0] finallayer_0_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_0_Im; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_1_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_1_Im; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_2_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_2_Im; // @[FFTDesigns.scala 421:31]
  FPComplexAdder FPComplexAdder ( // @[FFTDesigns.scala 258:34]
    .clock(FPComplexAdder_clock),
    .reset(FPComplexAdder_reset),
    .io_in_a_Re(FPComplexAdder_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_io_out_s_Im)
  );
  FPComplexSub FPComplexSub ( // @[FFTDesigns.scala 261:34]
    .clock(FPComplexSub_clock),
    .reset(FPComplexSub_reset),
    .io_in_a_Re(FPComplexSub_io_in_a_Re),
    .io_in_a_Im(FPComplexSub_io_in_a_Im),
    .io_in_b_Re(FPComplexSub_io_in_b_Re),
    .io_in_b_Im(FPComplexSub_io_in_b_Im),
    .io_out_s_Re(FPComplexSub_io_out_s_Re),
    .io_out_s_Im(FPComplexSub_io_out_s_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder ( // @[FFTDesigns.scala 275:36]
    .io_in_0_Re(FPComplexMultiAdder_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_io_out_Im)
  );
  FPComplexMult_reducable_v2 FPComplexMult_reducable_v2 ( // @[FFTDesigns.scala 294:39]
    .clock(FPComplexMult_reducable_v2_clock),
    .reset(FPComplexMult_reducable_v2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_1 FPComplexMult_reducable_v2_1 ( // @[FFTDesigns.scala 297:39]
    .clock(FPComplexMult_reducable_v2_1_clock),
    .reset(FPComplexMult_reducable_v2_1_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_1_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_1_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_reducable ( // @[FFTDesigns.scala 338:34]
    .clock(FPComplexAdder_reducable_clock),
    .reset(FPComplexAdder_reducable_reset),
    .io_in_a_Re(FPComplexAdder_reducable_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_reducable_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_reducable_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_reducable_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_reducable_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_reducable_io_out_s_Im)
  );
  FPComplexSub FPComplexSub_reducable ( // @[FFTDesigns.scala 341:34]
    .clock(FPComplexSub_reducable_clock),
    .reset(FPComplexSub_reducable_reset),
    .io_in_a_Re(FPComplexSub_reducable_io_in_a_Re),
    .io_in_a_Im(FPComplexSub_reducable_io_in_a_Im),
    .io_in_b_Re(FPComplexSub_reducable_io_in_b_Re),
    .io_in_b_Im(FPComplexSub_reducable_io_in_b_Im),
    .io_out_s_Re(FPComplexSub_reducable_io_out_s_Re),
    .io_out_s_Im(FPComplexSub_reducable_io_out_s_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder_1 ( // @[FFTDesigns.scala 394:29]
    .io_in_0_Re(FPComplexMultiAdder_1_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_1_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_1_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_1_io_out_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder_2 ( // @[FFTDesigns.scala 394:29]
    .io_in_0_Re(FPComplexMultiAdder_2_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_2_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_2_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_2_io_out_Im)
  );
  FPComplexAdder FPComplexAdder_1 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_1_clock),
    .reset(FPComplexAdder_1_reset),
    .io_in_a_Re(FPComplexAdder_1_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_1_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_1_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_1_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_1_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_1_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_2 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_2_clock),
    .reset(FPComplexAdder_2_reset),
    .io_in_a_Re(FPComplexAdder_2_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_2_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_2_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_2_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_2_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_2_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_3 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_3_clock),
    .reset(FPComplexAdder_3_reset),
    .io_in_a_Re(FPComplexAdder_3_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_3_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_3_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_3_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_3_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_3_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexAdder_1_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_0_Im = FPComplexAdder_1_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign io_out_1_Re = FPComplexAdder_2_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_1_Im = FPComplexAdder_2_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign io_out_2_Re = FPComplexAdder_3_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_2_Im = FPComplexAdder_3_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign FPComplexAdder_clock = clock;
  assign FPComplexAdder_reset = reset;
  assign FPComplexAdder_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 268:38]
  assign FPComplexAdder_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 268:38]
  assign FPComplexAdder_io_in_b_Re = io_in_2_Re; // @[FFTDesigns.scala 269:38]
  assign FPComplexAdder_io_in_b_Im = io_in_2_Im; // @[FFTDesigns.scala 269:38]
  assign FPComplexSub_clock = clock;
  assign FPComplexSub_reset = reset;
  assign FPComplexSub_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 270:38]
  assign FPComplexSub_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 270:38]
  assign FPComplexSub_io_in_b_Re = io_in_2_Re; // @[FFTDesigns.scala 271:38]
  assign FPComplexSub_io_in_b_Im = io_in_2_Im; // @[FFTDesigns.scala 271:38]
  assign FPComplexMultiAdder_io_in_0_Re = initial_layer_out_1_0_Re; // @[FFTDesigns.scala 290:27]
  assign FPComplexMultiAdder_io_in_0_Im = initial_layer_out_1_0_Im; // @[FFTDesigns.scala 290:27]
  assign FPComplexMult_reducable_v2_clock = clock;
  assign FPComplexMult_reducable_v2_reset = reset;
  assign FPComplexMult_reducable_v2_io_in_a_Re = FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 320:34]
  assign FPComplexMult_reducable_v2_io_in_a_Im = FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 320:34]
  assign FPComplexMult_reducable_v2_1_clock = clock;
  assign FPComplexMult_reducable_v2_1_reset = reset;
  assign FPComplexMult_reducable_v2_1_io_in_a_Re = FPComplexSub_io_out_s_Re; // @[FFTDesigns.scala 323:34]
  assign FPComplexMult_reducable_v2_1_io_in_a_Im = FPComplexSub_io_out_s_Im; // @[FFTDesigns.scala 323:34]
  assign FPComplexAdder_reducable_clock = clock;
  assign FPComplexAdder_reducable_reset = reset;
  assign FPComplexAdder_reducable_io_in_a_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 366:36]
  assign FPComplexAdder_reducable_io_in_a_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 366:36]
  assign FPComplexAdder_reducable_io_in_b_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 367:36]
  assign FPComplexAdder_reducable_io_in_b_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 367:36]
  assign FPComplexSub_reducable_clock = clock;
  assign FPComplexSub_reducable_reset = reset;
  assign FPComplexSub_reducable_io_in_a_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 368:36]
  assign FPComplexSub_reducable_io_in_a_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 368:36]
  assign FPComplexSub_reducable_io_in_b_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 369:36]
  assign FPComplexSub_reducable_io_in_b_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 369:36]
  assign FPComplexMultiAdder_1_io_in_0_Re = FPComplexAdder_reducable_io_out_s_Re; // @[FFTDesigns.scala 402:36]
  assign FPComplexMultiAdder_1_io_in_0_Im = FPComplexAdder_reducable_io_out_s_Im; // @[FFTDesigns.scala 402:36]
  assign FPComplexMultiAdder_2_io_in_0_Re = FPComplexSub_reducable_io_out_s_Re; // @[FFTDesigns.scala 404:61]
  assign FPComplexMultiAdder_2_io_in_0_Im = FPComplexSub_reducable_io_out_s_Im; // @[FFTDesigns.scala 404:61]
  assign FPComplexAdder_1_clock = clock;
  assign FPComplexAdder_1_reset = reset;
  assign FPComplexAdder_1_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_1_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_1_io_in_b_Re = FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_1_io_in_b_Im = FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_2_clock = clock;
  assign FPComplexAdder_2_reset = reset;
  assign FPComplexAdder_2_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_2_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_2_io_in_b_Re = FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_2_io_in_b_Im = FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_3_clock = clock;
  assign FPComplexAdder_3_reset = reset;
  assign FPComplexAdder_3_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_3_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_3_io_in_b_Re = FPComplexMultiAdder_2_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_3_io_in_b_Im = FPComplexMultiAdder_2_io_out_Im; // @[FFTDesigns.scala 431:35]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_0_0_Re <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_0_0_Re <= FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 281:37]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_0_0_Im <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_0_0_Im <= FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 281:37]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_1_0_Re <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_1_0_Re <= initial_layer_out_0_0_Re; // @[FFTDesigns.scala 284:32]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_1_0_Im <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_1_0_Im <= initial_layer_out_0_0_Im; // @[FFTDesigns.scala 284:32]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_0_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_0_Re <= io_in_0_Re; // @[FFTDesigns.scala 424:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_0_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_0_Im <= io_in_0_Im; // @[FFTDesigns.scala 424:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_1_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_1_Re <= finallayer_0_Re; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_1_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_1_Im <= finallayer_0_Im; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_2_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_2_Re <= finallayer_1_Re; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_2_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_2_Im <= finallayer_1_Im; // @[FFTDesigns.scala 426:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  initial_layer_out_0_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  initial_layer_out_0_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  initial_layer_out_1_0_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  initial_layer_out_1_0_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  finallayer_0_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  finallayer_0_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  finallayer_1_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  finallayer_1_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  finallayer_2_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  finallayer_2_Im = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PermutationsBasic(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im
);
  assign io_out_0_Re = io_in_0_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_0_Im = io_in_0_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Re = io_in_1_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Im = io_in_1_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Re = io_in_2_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Im = io_in_2_Im; // @[FFTDesigns.scala 2315:17]
endmodule
module FFT_sr_v2_nrv(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im
);
  wire  DFT_r_v2_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_2_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_2_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_2_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_2_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] PermutationsBasic_io_in_0_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_0_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_1_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_1_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_2_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_2_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_0_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_0_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_1_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_1_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_2_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_2_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_1_io_in_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_2_Im; // @[FFTDesigns.scala 3129:37]
  DFT_r_v2 DFT_r_v2 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_clock),
    .reset(DFT_r_v2_reset),
    .io_in_0_Re(DFT_r_v2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_io_out_2_Im)
  );
  PermutationsBasic PermutationsBasic ( // @[FFTDesigns.scala 3127:35]
    .io_in_0_Re(PermutationsBasic_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_io_in_2_Im),
    .io_out_0_Re(PermutationsBasic_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_io_out_2_Im)
  );
  PermutationsBasic PermutationsBasic_1 ( // @[FFTDesigns.scala 3129:37]
    .io_in_0_Re(PermutationsBasic_1_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_1_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_1_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_1_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_1_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_1_io_in_2_Im),
    .io_out_0_Re(PermutationsBasic_1_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_1_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_1_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_1_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_1_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_1_io_out_2_Im)
  );
  assign io_out_0_Re = PermutationsBasic_1_io_out_0_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_0_Im = PermutationsBasic_1_io_out_0_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_1_Re = PermutationsBasic_1_io_out_1_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_1_Im = PermutationsBasic_1_io_out_1_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_2_Re = PermutationsBasic_1_io_out_2_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_2_Im = PermutationsBasic_1_io_out_2_Im; // @[FFTDesigns.scala 3159:12]
  assign DFT_r_v2_clock = clock;
  assign DFT_r_v2_reset = reset;
  assign DFT_r_v2_io_in_0_Re = PermutationsBasic_io_out_0_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_io_in_0_Im = PermutationsBasic_io_out_0_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_io_in_1_Re = PermutationsBasic_io_out_1_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_io_in_1_Im = PermutationsBasic_io_out_1_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_io_in_2_Re = PermutationsBasic_io_out_2_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_io_in_2_Im = PermutationsBasic_io_out_2_Im; // @[FFTDesigns.scala 3145:39]
  assign PermutationsBasic_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_2_Re = io_in_2_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_2_Im = io_in_2_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_1_io_in_0_Re = DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_0_Im = DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_1_Re = DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_1_Im = DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_2_Re = DFT_r_v2_io_out_2_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_2_Im = DFT_r_v2_io_out_2_Im; // @[FFTDesigns.scala 3149:43]
endmodule
module FPComplexMultiAdder_96(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  wire  FPComplexAdder_clock; // @[FPComplex.scala 477:30]
  wire  FPComplexAdder_reset; // @[FPComplex.scala 477:30]
  wire [31:0] FPComplexAdder_io_in_a_Re; // @[FPComplex.scala 477:30]
  wire [31:0] FPComplexAdder_io_in_a_Im; // @[FPComplex.scala 477:30]
  wire [31:0] FPComplexAdder_io_in_b_Re; // @[FPComplex.scala 477:30]
  wire [31:0] FPComplexAdder_io_in_b_Im; // @[FPComplex.scala 477:30]
  wire [31:0] FPComplexAdder_io_out_s_Re; // @[FPComplex.scala 477:30]
  wire [31:0] FPComplexAdder_io_out_s_Im; // @[FPComplex.scala 477:30]
  FPComplexAdder FPComplexAdder ( // @[FPComplex.scala 477:30]
    .clock(FPComplexAdder_clock),
    .reset(FPComplexAdder_reset),
    .io_in_a_Re(FPComplexAdder_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_io_out_s_Im)
  );
  assign io_out_Re = FPComplexAdder_io_out_s_Re; // @[FPComplex.scala 595:16]
  assign io_out_Im = FPComplexAdder_io_out_s_Im; // @[FPComplex.scala 595:16]
  assign FPComplexAdder_clock = clock;
  assign FPComplexAdder_reset = reset;
  assign FPComplexAdder_io_in_a_Re = io_in_0_Re; // @[FPComplex.scala 557:42]
  assign FPComplexAdder_io_in_a_Im = io_in_0_Im; // @[FPComplex.scala 557:42]
  assign FPComplexAdder_io_in_b_Re = io_in_1_Re; // @[FPComplex.scala 558:42]
  assign FPComplexAdder_io_in_b_Im = io_in_1_Im; // @[FPComplex.scala 558:42]
endmodule
module DFT_r_V1_nonregout(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im
);
  wire [31:0] cmplx_adj_io_in_Re; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_in_Im; // @[FFTDesigns.scala 1808:22]
  wire [7:0] cmplx_adj_io_in_adj; // @[FFTDesigns.scala 1808:22]
  wire  cmplx_adj_io_is_neg; // @[FFTDesigns.scala 1808:22]
  wire  cmplx_adj_io_is_flip; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_out_Re; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_out_Im; // @[FFTDesigns.scala 1808:22]
  wire  FPComplexMultiAdder_clock; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_reset; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_0_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_0_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_1_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_1_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_1_clock; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_1_reset; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_1_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_1_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 1839:26]
  cmplx_adj cmplx_adj ( // @[FFTDesigns.scala 1808:22]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  FPComplexMultiAdder_96 FPComplexMultiAdder ( // @[FFTDesigns.scala 1839:26]
    .clock(FPComplexMultiAdder_clock),
    .reset(FPComplexMultiAdder_reset),
    .io_in_0_Re(FPComplexMultiAdder_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_io_in_1_Im),
    .io_out_Re(FPComplexMultiAdder_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_io_out_Im)
  );
  FPComplexMultiAdder_96 FPComplexMultiAdder_1 ( // @[FFTDesigns.scala 1839:26]
    .clock(FPComplexMultiAdder_1_clock),
    .reset(FPComplexMultiAdder_1_reset),
    .io_in_0_Re(FPComplexMultiAdder_1_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_1_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_1_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_1_io_in_1_Im),
    .io_out_Re(FPComplexMultiAdder_1_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_1_io_out_Im)
  );
  assign io_out_0_Re = FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 1911:17]
  assign io_out_0_Im = FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 1911:17]
  assign io_out_1_Re = FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 1911:17]
  assign io_out_1_Im = FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 1911:17]
  assign cmplx_adj_io_in_Re = io_in_1_Re; // @[FFTDesigns.scala 1820:27]
  assign cmplx_adj_io_in_Im = io_in_1_Im; // @[FFTDesigns.scala 1820:27]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FFTDesigns.scala 1821:31]
  assign cmplx_adj_io_is_neg = 1'h1; // @[FFTDesigns.scala 1822:31]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FFTDesigns.scala 1823:32]
  assign FPComplexMultiAdder_clock = clock;
  assign FPComplexMultiAdder_reset = reset;
  assign FPComplexMultiAdder_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_1_clock = clock;
  assign FPComplexMultiAdder_1_reset = reset;
  assign FPComplexMultiAdder_1_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 1896:32]
  assign FPComplexMultiAdder_1_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 1896:32]
  assign FPComplexMultiAdder_1_io_in_1_Re = cmplx_adj_io_out_Re; // @[FFTDesigns.scala 1818:24 1824:42]
  assign FPComplexMultiAdder_1_io_in_1_Im = cmplx_adj_io_out_Im; // @[FFTDesigns.scala 1818:24 1824:42]
endmodule
module DFT_r_v2_32(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im
);
  wire  DFT_r_V1_nonregout_clock; // @[FFTDesigns.scala 169:24]
  wire  DFT_r_V1_nonregout_reset; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_0_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_0_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_1_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_1_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_0_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_0_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_1_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_1_Im; // @[FFTDesigns.scala 169:24]
  DFT_r_V1_nonregout DFT_r_V1_nonregout ( // @[FFTDesigns.scala 169:24]
    .clock(DFT_r_V1_nonregout_clock),
    .reset(DFT_r_V1_nonregout_reset),
    .io_in_0_Re(DFT_r_V1_nonregout_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_nonregout_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_nonregout_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_nonregout_io_in_1_Im),
    .io_out_0_Re(DFT_r_V1_nonregout_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_nonregout_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_nonregout_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_nonregout_io_out_1_Im)
  );
  assign io_out_0_Re = DFT_r_V1_nonregout_io_out_0_Re; // @[FFTDesigns.scala 171:14]
  assign io_out_0_Im = DFT_r_V1_nonregout_io_out_0_Im; // @[FFTDesigns.scala 171:14]
  assign io_out_1_Re = DFT_r_V1_nonregout_io_out_1_Re; // @[FFTDesigns.scala 171:14]
  assign io_out_1_Im = DFT_r_V1_nonregout_io_out_1_Im; // @[FFTDesigns.scala 171:14]
  assign DFT_r_V1_nonregout_clock = clock;
  assign DFT_r_V1_nonregout_reset = reset;
  assign DFT_r_V1_nonregout_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 170:15]
endmodule
module PermutationsBasic_64(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im
);
  assign io_out_0_Re = io_in_0_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_0_Im = io_in_0_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Re = io_in_16_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Im = io_in_16_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Re = io_in_8_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Im = io_in_8_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_3_Re = io_in_24_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_3_Im = io_in_24_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_4_Re = io_in_4_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_4_Im = io_in_4_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_5_Re = io_in_20_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_5_Im = io_in_20_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_6_Re = io_in_12_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_6_Im = io_in_12_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_7_Re = io_in_28_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_7_Im = io_in_28_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_8_Re = io_in_2_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_8_Im = io_in_2_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_9_Re = io_in_18_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_9_Im = io_in_18_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_10_Re = io_in_10_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_10_Im = io_in_10_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_11_Re = io_in_26_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_11_Im = io_in_26_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_12_Re = io_in_6_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_12_Im = io_in_6_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_13_Re = io_in_22_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_13_Im = io_in_22_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_14_Re = io_in_14_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_14_Im = io_in_14_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_15_Re = io_in_30_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_15_Im = io_in_30_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_16_Re = io_in_1_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_16_Im = io_in_1_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_17_Re = io_in_17_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_17_Im = io_in_17_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_18_Re = io_in_9_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_18_Im = io_in_9_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_19_Re = io_in_25_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_19_Im = io_in_25_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_20_Re = io_in_5_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_20_Im = io_in_5_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_21_Re = io_in_21_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_21_Im = io_in_21_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_22_Re = io_in_13_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_22_Im = io_in_13_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_23_Re = io_in_29_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_23_Im = io_in_29_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_24_Re = io_in_3_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_24_Im = io_in_3_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_25_Re = io_in_19_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_25_Im = io_in_19_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_26_Re = io_in_11_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_26_Im = io_in_11_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_27_Re = io_in_27_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_27_Im = io_in_27_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_28_Re = io_in_7_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_28_Im = io_in_7_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_29_Re = io_in_23_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_29_Im = io_in_23_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_30_Re = io_in_15_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_30_Im = io_in_15_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_31_Re = io_in_31_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_31_Im = io_in_31_Im; // @[FFTDesigns.scala 2315:17]
endmodule
module PermutationsBasic_65(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im
);
  assign io_out_0_Re = io_in_0_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_0_Im = io_in_0_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Re = io_in_2_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Im = io_in_2_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Re = io_in_4_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Im = io_in_4_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_3_Re = io_in_6_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_3_Im = io_in_6_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_4_Re = io_in_8_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_4_Im = io_in_8_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_5_Re = io_in_10_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_5_Im = io_in_10_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_6_Re = io_in_12_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_6_Im = io_in_12_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_7_Re = io_in_14_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_7_Im = io_in_14_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_8_Re = io_in_16_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_8_Im = io_in_16_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_9_Re = io_in_18_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_9_Im = io_in_18_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_10_Re = io_in_20_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_10_Im = io_in_20_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_11_Re = io_in_22_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_11_Im = io_in_22_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_12_Re = io_in_24_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_12_Im = io_in_24_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_13_Re = io_in_26_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_13_Im = io_in_26_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_14_Re = io_in_28_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_14_Im = io_in_28_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_15_Re = io_in_30_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_15_Im = io_in_30_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_16_Re = io_in_1_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_16_Im = io_in_1_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_17_Re = io_in_3_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_17_Im = io_in_3_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_18_Re = io_in_5_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_18_Im = io_in_5_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_19_Re = io_in_7_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_19_Im = io_in_7_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_20_Re = io_in_9_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_20_Im = io_in_9_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_21_Re = io_in_11_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_21_Im = io_in_11_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_22_Re = io_in_13_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_22_Im = io_in_13_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_23_Re = io_in_15_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_23_Im = io_in_15_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_24_Re = io_in_17_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_24_Im = io_in_17_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_25_Re = io_in_19_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_25_Im = io_in_19_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_26_Re = io_in_21_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_26_Im = io_in_21_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_27_Re = io_in_23_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_27_Im = io_in_23_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_28_Re = io_in_25_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_28_Im = io_in_25_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_29_Re = io_in_27_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_29_Im = io_in_27_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_30_Re = io_in_29_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_30_Im = io_in_29_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_31_Re = io_in_31_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_31_Im = io_in_31_Im; // @[FFTDesigns.scala 2315:17]
endmodule
module FPComplexMult_reducable_v2_64(
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 333:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 333:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 333:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 333:33]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 333:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  assign io_out_s_Re = cmplx_adj_io_out_Re; // @[FPComplex.scala 355:20]
  assign io_out_s_Im = cmplx_adj_io_out_Im; // @[FPComplex.scala 355:20]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 334:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 334:24]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FPComplex.scala 337:30]
  assign cmplx_adj_io_is_neg = 1'h0; // @[FPComplex.scala 341:32]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FPComplex.scala 335:29]
endmodule
module FPComplexMult_reducable_v2_81(
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 293:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 293:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 293:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 293:33]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 293:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  assign io_out_s_Re = cmplx_adj_io_out_Re; // @[FPComplex.scala 315:20]
  assign io_out_s_Im = cmplx_adj_io_out_Im; // @[FPComplex.scala 315:20]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 294:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 294:24]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FPComplex.scala 297:30]
  assign cmplx_adj_io_is_neg = 1'h1; // @[FPComplex.scala 299:32]
  assign cmplx_adj_io_is_flip = 1'h1; // @[FPComplex.scala 295:29]
endmodule
module TwiddleFactors(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im
);
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_1 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_1_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_1_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_2 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_3 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_3_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_3_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_4 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_4_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_4_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_5 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_5_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_5_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_6 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_6_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_6_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_7 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_7_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_7_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_8 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_8_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_8_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_9 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_9_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_9_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_10 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_10_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_10_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_11 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_11_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_11_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_12 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_12_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_12_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_13 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_13_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_13_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_14 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_14_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_14_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_15 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_15_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_15_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_16 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_16_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_16_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_16_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_16_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_81 FPComplexMult_reducable_v2_17 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_17_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_17_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_17_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_17_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_18 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_18_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_18_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_18_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_18_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_81 FPComplexMult_reducable_v2_19 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_19_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_19_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_19_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_19_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_20 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_20_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_20_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_20_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_20_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_81 FPComplexMult_reducable_v2_21 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_21_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_21_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_21_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_21_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_22 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_22_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_22_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_22_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_22_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_81 FPComplexMult_reducable_v2_23 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_23_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_23_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_23_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_23_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_24 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_24_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_24_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_24_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_24_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_81 FPComplexMult_reducable_v2_25 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_25_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_25_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_25_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_25_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_26 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_26_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_26_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_26_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_26_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_81 FPComplexMult_reducable_v2_27 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_27_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_27_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_27_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_27_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_28 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_28_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_28_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_28_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_28_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_81 FPComplexMult_reducable_v2_29 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_29_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_29_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_29_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_29_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_64 FPComplexMult_reducable_v2_30 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_30_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_30_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_30_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_30_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_81 FPComplexMult_reducable_v2_31 ( // @[FFTDesigns.scala 2298:28]
    .io_in_a_Re(FPComplexMult_reducable_v2_31_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_31_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_31_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_31_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_0_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_1_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_1_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_2_Re = FPComplexMult_reducable_v2_2_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_2_Im = FPComplexMult_reducable_v2_2_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_3_Re = FPComplexMult_reducable_v2_3_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_3_Im = FPComplexMult_reducable_v2_3_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_4_Re = FPComplexMult_reducable_v2_4_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_4_Im = FPComplexMult_reducable_v2_4_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_5_Re = FPComplexMult_reducable_v2_5_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_5_Im = FPComplexMult_reducable_v2_5_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_6_Re = FPComplexMult_reducable_v2_6_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_6_Im = FPComplexMult_reducable_v2_6_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_7_Re = FPComplexMult_reducable_v2_7_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_7_Im = FPComplexMult_reducable_v2_7_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_8_Re = FPComplexMult_reducable_v2_8_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_8_Im = FPComplexMult_reducable_v2_8_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_9_Re = FPComplexMult_reducable_v2_9_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_9_Im = FPComplexMult_reducable_v2_9_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_10_Re = FPComplexMult_reducable_v2_10_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_10_Im = FPComplexMult_reducable_v2_10_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_11_Re = FPComplexMult_reducable_v2_11_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_11_Im = FPComplexMult_reducable_v2_11_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_12_Re = FPComplexMult_reducable_v2_12_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_12_Im = FPComplexMult_reducable_v2_12_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_13_Re = FPComplexMult_reducable_v2_13_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_13_Im = FPComplexMult_reducable_v2_13_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_14_Re = FPComplexMult_reducable_v2_14_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_14_Im = FPComplexMult_reducable_v2_14_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_15_Re = FPComplexMult_reducable_v2_15_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_15_Im = FPComplexMult_reducable_v2_15_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_16_Re = FPComplexMult_reducable_v2_16_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_16_Im = FPComplexMult_reducable_v2_16_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_17_Re = FPComplexMult_reducable_v2_17_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_17_Im = FPComplexMult_reducable_v2_17_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_18_Re = FPComplexMult_reducable_v2_18_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_18_Im = FPComplexMult_reducable_v2_18_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_19_Re = FPComplexMult_reducable_v2_19_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_19_Im = FPComplexMult_reducable_v2_19_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_20_Re = FPComplexMult_reducable_v2_20_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_20_Im = FPComplexMult_reducable_v2_20_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_21_Re = FPComplexMult_reducable_v2_21_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_21_Im = FPComplexMult_reducable_v2_21_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_22_Re = FPComplexMult_reducable_v2_22_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_22_Im = FPComplexMult_reducable_v2_22_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_23_Re = FPComplexMult_reducable_v2_23_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_23_Im = FPComplexMult_reducable_v2_23_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_24_Re = FPComplexMult_reducable_v2_24_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_24_Im = FPComplexMult_reducable_v2_24_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_25_Re = FPComplexMult_reducable_v2_25_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_25_Im = FPComplexMult_reducable_v2_25_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_26_Re = FPComplexMult_reducable_v2_26_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_26_Im = FPComplexMult_reducable_v2_26_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_27_Re = FPComplexMult_reducable_v2_27_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_27_Im = FPComplexMult_reducable_v2_27_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_28_Re = FPComplexMult_reducable_v2_28_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_28_Im = FPComplexMult_reducable_v2_28_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_29_Re = FPComplexMult_reducable_v2_29_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_29_Im = FPComplexMult_reducable_v2_29_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_30_Re = FPComplexMult_reducable_v2_30_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_30_Im = FPComplexMult_reducable_v2_30_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_31_Re = FPComplexMult_reducable_v2_31_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_31_Im = FPComplexMult_reducable_v2_31_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign FPComplexMult_reducable_v2_io_in_a_Re = io_in_0_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_io_in_a_Im = io_in_0_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_1_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_1_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_2_io_in_a_Re = io_in_2_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_2_io_in_a_Im = io_in_2_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_io_in_a_Re = io_in_3_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_io_in_a_Im = io_in_3_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_4_io_in_a_Re = io_in_4_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_4_io_in_a_Im = io_in_4_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_io_in_a_Re = io_in_5_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_io_in_a_Im = io_in_5_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_6_io_in_a_Re = io_in_6_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_6_io_in_a_Im = io_in_6_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_io_in_a_Re = io_in_7_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_io_in_a_Im = io_in_7_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_8_io_in_a_Re = io_in_8_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_8_io_in_a_Im = io_in_8_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_io_in_a_Re = io_in_9_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_io_in_a_Im = io_in_9_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_10_io_in_a_Re = io_in_10_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_10_io_in_a_Im = io_in_10_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_io_in_a_Re = io_in_11_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_io_in_a_Im = io_in_11_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_12_io_in_a_Re = io_in_12_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_12_io_in_a_Im = io_in_12_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_io_in_a_Re = io_in_13_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_io_in_a_Im = io_in_13_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_14_io_in_a_Re = io_in_14_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_14_io_in_a_Im = io_in_14_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_io_in_a_Re = io_in_15_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_io_in_a_Im = io_in_15_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_16_io_in_a_Re = io_in_16_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_16_io_in_a_Im = io_in_16_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_17_io_in_a_Re = io_in_17_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_17_io_in_a_Im = io_in_17_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_18_io_in_a_Re = io_in_18_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_18_io_in_a_Im = io_in_18_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_io_in_a_Re = io_in_19_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_io_in_a_Im = io_in_19_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_20_io_in_a_Re = io_in_20_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_20_io_in_a_Im = io_in_20_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_io_in_a_Re = io_in_21_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_io_in_a_Im = io_in_21_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_22_io_in_a_Re = io_in_22_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_22_io_in_a_Im = io_in_22_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_io_in_a_Re = io_in_23_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_io_in_a_Im = io_in_23_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_24_io_in_a_Re = io_in_24_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_24_io_in_a_Im = io_in_24_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_io_in_a_Re = io_in_25_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_io_in_a_Im = io_in_25_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_26_io_in_a_Re = io_in_26_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_26_io_in_a_Im = io_in_26_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_io_in_a_Re = io_in_27_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_io_in_a_Im = io_in_27_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_28_io_in_a_Re = io_in_28_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_28_io_in_a_Im = io_in_28_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_io_in_a_Re = io_in_29_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_io_in_a_Im = io_in_29_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_30_io_in_a_Re = io_in_30_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_30_io_in_a_Im = io_in_30_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_io_in_a_Re = io_in_31_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_io_in_a_Im = io_in_31_Im; // @[FFTDesigns.scala 2302:27]
endmodule
module FPComplexMult_reducable_v2_96(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 333:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 333:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 333:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 333:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 333:33]
  reg [31:0] result_0_Re; // @[FPComplex.scala 344:31]
  reg [31:0] result_0_Im; // @[FPComplex.scala 344:31]
  reg [31:0] result_1_Re; // @[FPComplex.scala 344:31]
  reg [31:0] result_1_Im; // @[FPComplex.scala 344:31]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 333:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  assign io_out_s_Re = result_1_Re; // @[FPComplex.scala 353:20]
  assign io_out_s_Im = result_1_Im; // @[FPComplex.scala 353:20]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 334:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 334:24]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FPComplex.scala 337:30]
  assign cmplx_adj_io_is_neg = 1'h0; // @[FPComplex.scala 341:32]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FPComplex.scala 335:29]
  always @(posedge clock) begin
    if (reset) begin // @[FPComplex.scala 344:31]
      result_0_Re <= 32'h0; // @[FPComplex.scala 344:31]
    end else begin
      result_0_Re <= cmplx_adj_io_out_Re; // @[FPComplex.scala 347:25]
    end
    if (reset) begin // @[FPComplex.scala 344:31]
      result_0_Im <= 32'h0; // @[FPComplex.scala 344:31]
    end else begin
      result_0_Im <= cmplx_adj_io_out_Im; // @[FPComplex.scala 347:25]
    end
    if (reset) begin // @[FPComplex.scala 344:31]
      result_1_Re <= 32'h0; // @[FPComplex.scala 344:31]
    end else begin
      result_1_Re <= result_0_Re; // @[FPComplex.scala 349:25]
    end
    if (reset) begin // @[FPComplex.scala 344:31]
      result_1_Im <= 32'h0; // @[FPComplex.scala 344:31]
    end else begin
      result_1_Im <= result_0_Im; // @[FPComplex.scala 349:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  result_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  result_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  result_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  result_1_Im = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMult_reducable_v2_105(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_subber_clock; // @[FPComplex.scala 372:26]
  wire  FP_subber_reset; // @[FPComplex.scala 372:26]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 372:26]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 372:26]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 372:26]
  wire  FP_adder_clock; // @[FPComplex.scala 373:26]
  wire  FP_adder_reset; // @[FPComplex.scala 373:26]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 373:26]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 373:26]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 373:26]
  wire  FP_multiplier_clock; // @[FPComplex.scala 431:30]
  wire  FP_multiplier_reset; // @[FPComplex.scala 431:30]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 431:30]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 431:30]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 431:30]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 431:30]
  wire  FP_multiplier_1_reset; // @[FPComplex.scala 431:30]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 431:30]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 431:30]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 431:30]
  wire  FP_multiplier_2_clock; // @[FPComplex.scala 450:30]
  wire  FP_multiplier_2_reset; // @[FPComplex.scala 450:30]
  wire [31:0] FP_multiplier_2_io_in_a; // @[FPComplex.scala 450:30]
  wire [31:0] FP_multiplier_2_io_in_b; // @[FPComplex.scala 450:30]
  wire [31:0] FP_multiplier_2_io_out_s; // @[FPComplex.scala 450:30]
  wire  FP_multiplier_3_clock; // @[FPComplex.scala 450:30]
  wire  FP_multiplier_3_reset; // @[FPComplex.scala 450:30]
  wire [31:0] FP_multiplier_3_io_in_a; // @[FPComplex.scala 450:30]
  wire [31:0] FP_multiplier_3_io_in_b; // @[FPComplex.scala 450:30]
  wire [31:0] FP_multiplier_3_io_out_s; // @[FPComplex.scala 450:30]
  FP_subber FP_subber ( // @[FPComplex.scala 372:26]
    .clock(FP_subber_clock),
    .reset(FP_subber_reset),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_adder FP_adder ( // @[FPComplex.scala 373:26]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 431:30]
    .clock(FP_multiplier_clock),
    .reset(FP_multiplier_reset),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 431:30]
    .clock(FP_multiplier_1_clock),
    .reset(FP_multiplier_1_reset),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  FP_multiplier FP_multiplier_2 ( // @[FPComplex.scala 450:30]
    .clock(FP_multiplier_2_clock),
    .reset(FP_multiplier_2_reset),
    .io_in_a(FP_multiplier_2_io_in_a),
    .io_in_b(FP_multiplier_2_io_in_b),
    .io_out_s(FP_multiplier_2_io_out_s)
  );
  FP_multiplier FP_multiplier_3 ( // @[FPComplex.scala 450:30]
    .clock(FP_multiplier_3_clock),
    .reset(FP_multiplier_3_reset),
    .io_in_a(FP_multiplier_3_io_in_a),
    .io_in_b(FP_multiplier_3_io_in_b),
    .io_out_s(FP_multiplier_3_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 464:19]
  assign io_out_s_Im = FP_adder_io_out_s; // @[FPComplex.scala 465:19]
  assign FP_subber_clock = clock;
  assign FP_subber_reset = reset;
  assign FP_subber_io_in_a = FP_multiplier_io_out_s; // @[FPComplex.scala 421:30 438:25]
  assign FP_subber_io_in_b = FP_multiplier_3_io_out_s; // @[FPComplex.scala 421:30 458:25]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = FP_multiplier_2_io_out_s; // @[FPComplex.scala 421:30 457:25]
  assign FP_adder_io_in_b = FP_multiplier_1_io_out_s; // @[FPComplex.scala 421:30 439:25]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_reset = reset;
  assign FP_multiplier_io_in_a = io_in_a_Re; // @[FPComplex.scala 434:33]
  assign FP_multiplier_io_in_b = io_in_b_Re; // @[FPComplex.scala 435:33]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_reset = reset;
  assign FP_multiplier_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 436:33]
  assign FP_multiplier_1_io_in_b = io_in_b_Re; // @[FPComplex.scala 437:33]
  assign FP_multiplier_2_clock = clock;
  assign FP_multiplier_2_reset = reset;
  assign FP_multiplier_2_io_in_a = io_in_a_Re; // @[FPComplex.scala 453:33]
  assign FP_multiplier_2_io_in_b = io_in_b_Im; // @[FPComplex.scala 454:33]
  assign FP_multiplier_3_clock = clock;
  assign FP_multiplier_3_reset = reset;
  assign FP_multiplier_3_io_in_a = io_in_a_Im; // @[FPComplex.scala 455:33]
  assign FP_multiplier_3_io_in_b = io_in_b_Im; // @[FPComplex.scala 456:33]
endmodule
module FPComplexMult_reducable_v2_113(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 293:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 293:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 293:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 293:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 293:33]
  reg [31:0] result_0_Re; // @[FPComplex.scala 304:31]
  reg [31:0] result_0_Im; // @[FPComplex.scala 304:31]
  reg [31:0] result_1_Re; // @[FPComplex.scala 304:31]
  reg [31:0] result_1_Im; // @[FPComplex.scala 304:31]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 293:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  assign io_out_s_Re = result_1_Re; // @[FPComplex.scala 313:20]
  assign io_out_s_Im = result_1_Im; // @[FPComplex.scala 313:20]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 294:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 294:24]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FPComplex.scala 297:30]
  assign cmplx_adj_io_is_neg = 1'h1; // @[FPComplex.scala 299:32]
  assign cmplx_adj_io_is_flip = 1'h1; // @[FPComplex.scala 295:29]
  always @(posedge clock) begin
    if (reset) begin // @[FPComplex.scala 304:31]
      result_0_Re <= 32'h0; // @[FPComplex.scala 304:31]
    end else begin
      result_0_Re <= cmplx_adj_io_out_Re; // @[FPComplex.scala 307:25]
    end
    if (reset) begin // @[FPComplex.scala 304:31]
      result_0_Im <= 32'h0; // @[FPComplex.scala 304:31]
    end else begin
      result_0_Im <= cmplx_adj_io_out_Im; // @[FPComplex.scala 307:25]
    end
    if (reset) begin // @[FPComplex.scala 304:31]
      result_1_Re <= 32'h0; // @[FPComplex.scala 304:31]
    end else begin
      result_1_Re <= result_0_Re; // @[FPComplex.scala 309:25]
    end
    if (reset) begin // @[FPComplex.scala 304:31]
      result_1_Im <= 32'h0; // @[FPComplex.scala 304:31]
    end else begin
      result_1_Im <= result_0_Im; // @[FPComplex.scala 309:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  result_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  result_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  result_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  result_1_Im = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactors_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im
);
  wire  FPComplexMult_reducable_v2_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_1_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_1_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_2_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_2_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_3_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_3_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_4_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_4_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_5_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_5_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_6_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_6_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_7_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_7_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_8_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_8_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_9_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_9_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_10_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_10_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_11_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_11_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_12_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_12_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_13_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_13_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_14_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_14_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_15_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_15_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_16_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_16_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_17_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_17_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_18_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_18_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_19_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_19_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_20_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_20_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_21_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_21_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_22_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_22_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_23_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_23_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_24_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_24_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_25_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_25_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_26_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_26_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_27_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_27_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_28_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_28_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_29_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_29_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_30_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_30_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_31_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_31_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_clock),
    .reset(FPComplexMult_reducable_v2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_1 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_1_clock),
    .reset(FPComplexMult_reducable_v2_1_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_1_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_1_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_2 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_2_clock),
    .reset(FPComplexMult_reducable_v2_2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_3 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_3_clock),
    .reset(FPComplexMult_reducable_v2_3_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_3_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_3_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_4 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_4_clock),
    .reset(FPComplexMult_reducable_v2_4_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_4_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_4_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_5 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_5_clock),
    .reset(FPComplexMult_reducable_v2_5_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_5_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_5_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_6 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_6_clock),
    .reset(FPComplexMult_reducable_v2_6_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_6_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_6_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_7 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_7_clock),
    .reset(FPComplexMult_reducable_v2_7_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_7_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_7_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_8 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_8_clock),
    .reset(FPComplexMult_reducable_v2_8_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_8_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_8_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_9 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_9_clock),
    .reset(FPComplexMult_reducable_v2_9_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_9_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_10 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_10_clock),
    .reset(FPComplexMult_reducable_v2_10_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_10_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_10_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_11 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_11_clock),
    .reset(FPComplexMult_reducable_v2_11_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_11_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_12 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_12_clock),
    .reset(FPComplexMult_reducable_v2_12_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_12_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_12_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_13 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_13_clock),
    .reset(FPComplexMult_reducable_v2_13_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_13_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_14 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_14_clock),
    .reset(FPComplexMult_reducable_v2_14_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_14_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_14_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_15 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_15_clock),
    .reset(FPComplexMult_reducable_v2_15_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_15_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_16 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_16_clock),
    .reset(FPComplexMult_reducable_v2_16_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_16_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_16_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_16_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_16_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_113 FPComplexMult_reducable_v2_17 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_17_clock),
    .reset(FPComplexMult_reducable_v2_17_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_17_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_17_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_17_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_17_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_18 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_18_clock),
    .reset(FPComplexMult_reducable_v2_18_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_18_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_18_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_18_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_18_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_113 FPComplexMult_reducable_v2_19 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_19_clock),
    .reset(FPComplexMult_reducable_v2_19_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_19_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_19_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_19_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_19_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_20 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_20_clock),
    .reset(FPComplexMult_reducable_v2_20_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_20_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_20_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_20_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_20_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_113 FPComplexMult_reducable_v2_21 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_21_clock),
    .reset(FPComplexMult_reducable_v2_21_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_21_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_21_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_21_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_21_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_22 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_22_clock),
    .reset(FPComplexMult_reducable_v2_22_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_22_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_22_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_22_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_22_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_113 FPComplexMult_reducable_v2_23 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_23_clock),
    .reset(FPComplexMult_reducable_v2_23_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_23_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_23_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_23_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_23_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_24 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_24_clock),
    .reset(FPComplexMult_reducable_v2_24_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_24_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_24_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_24_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_24_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_25 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_25_clock),
    .reset(FPComplexMult_reducable_v2_25_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_25_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_25_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_25_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_25_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_25_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_25_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_26 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_26_clock),
    .reset(FPComplexMult_reducable_v2_26_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_26_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_26_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_26_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_26_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_27 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_27_clock),
    .reset(FPComplexMult_reducable_v2_27_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_27_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_27_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_27_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_27_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_27_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_27_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_28 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_28_clock),
    .reset(FPComplexMult_reducable_v2_28_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_28_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_28_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_28_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_28_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_29 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_29_clock),
    .reset(FPComplexMult_reducable_v2_29_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_29_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_29_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_29_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_29_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_29_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_29_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_30 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_30_clock),
    .reset(FPComplexMult_reducable_v2_30_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_30_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_30_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_30_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_30_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_31 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_31_clock),
    .reset(FPComplexMult_reducable_v2_31_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_31_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_31_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_31_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_31_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_31_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_31_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_0_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_1_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_1_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_2_Re = FPComplexMult_reducable_v2_2_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_2_Im = FPComplexMult_reducable_v2_2_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_3_Re = FPComplexMult_reducable_v2_3_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_3_Im = FPComplexMult_reducable_v2_3_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_4_Re = FPComplexMult_reducable_v2_4_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_4_Im = FPComplexMult_reducable_v2_4_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_5_Re = FPComplexMult_reducable_v2_5_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_5_Im = FPComplexMult_reducable_v2_5_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_6_Re = FPComplexMult_reducable_v2_6_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_6_Im = FPComplexMult_reducable_v2_6_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_7_Re = FPComplexMult_reducable_v2_7_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_7_Im = FPComplexMult_reducable_v2_7_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_8_Re = FPComplexMult_reducable_v2_8_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_8_Im = FPComplexMult_reducable_v2_8_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_9_Re = FPComplexMult_reducable_v2_9_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_9_Im = FPComplexMult_reducable_v2_9_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_10_Re = FPComplexMult_reducable_v2_10_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_10_Im = FPComplexMult_reducable_v2_10_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_11_Re = FPComplexMult_reducable_v2_11_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_11_Im = FPComplexMult_reducable_v2_11_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_12_Re = FPComplexMult_reducable_v2_12_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_12_Im = FPComplexMult_reducable_v2_12_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_13_Re = FPComplexMult_reducable_v2_13_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_13_Im = FPComplexMult_reducable_v2_13_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_14_Re = FPComplexMult_reducable_v2_14_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_14_Im = FPComplexMult_reducable_v2_14_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_15_Re = FPComplexMult_reducable_v2_15_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_15_Im = FPComplexMult_reducable_v2_15_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_16_Re = FPComplexMult_reducable_v2_16_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_16_Im = FPComplexMult_reducable_v2_16_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_17_Re = FPComplexMult_reducable_v2_17_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_17_Im = FPComplexMult_reducable_v2_17_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_18_Re = FPComplexMult_reducable_v2_18_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_18_Im = FPComplexMult_reducable_v2_18_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_19_Re = FPComplexMult_reducable_v2_19_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_19_Im = FPComplexMult_reducable_v2_19_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_20_Re = FPComplexMult_reducable_v2_20_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_20_Im = FPComplexMult_reducable_v2_20_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_21_Re = FPComplexMult_reducable_v2_21_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_21_Im = FPComplexMult_reducable_v2_21_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_22_Re = FPComplexMult_reducable_v2_22_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_22_Im = FPComplexMult_reducable_v2_22_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_23_Re = FPComplexMult_reducable_v2_23_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_23_Im = FPComplexMult_reducable_v2_23_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_24_Re = FPComplexMult_reducable_v2_24_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_24_Im = FPComplexMult_reducable_v2_24_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_25_Re = FPComplexMult_reducable_v2_25_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_25_Im = FPComplexMult_reducable_v2_25_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_26_Re = FPComplexMult_reducable_v2_26_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_26_Im = FPComplexMult_reducable_v2_26_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_27_Re = FPComplexMult_reducable_v2_27_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_27_Im = FPComplexMult_reducable_v2_27_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_28_Re = FPComplexMult_reducable_v2_28_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_28_Im = FPComplexMult_reducable_v2_28_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_29_Re = FPComplexMult_reducable_v2_29_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_29_Im = FPComplexMult_reducable_v2_29_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_30_Re = FPComplexMult_reducable_v2_30_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_30_Im = FPComplexMult_reducable_v2_30_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_31_Re = FPComplexMult_reducable_v2_31_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_31_Im = FPComplexMult_reducable_v2_31_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign FPComplexMult_reducable_v2_clock = clock;
  assign FPComplexMult_reducable_v2_reset = reset;
  assign FPComplexMult_reducable_v2_io_in_a_Re = io_in_0_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_io_in_a_Im = io_in_0_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_1_clock = clock;
  assign FPComplexMult_reducable_v2_1_reset = reset;
  assign FPComplexMult_reducable_v2_1_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_1_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_2_clock = clock;
  assign FPComplexMult_reducable_v2_2_reset = reset;
  assign FPComplexMult_reducable_v2_2_io_in_a_Re = io_in_2_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_2_io_in_a_Im = io_in_2_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_clock = clock;
  assign FPComplexMult_reducable_v2_3_reset = reset;
  assign FPComplexMult_reducable_v2_3_io_in_a_Re = io_in_3_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_io_in_a_Im = io_in_3_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_4_clock = clock;
  assign FPComplexMult_reducable_v2_4_reset = reset;
  assign FPComplexMult_reducable_v2_4_io_in_a_Re = io_in_4_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_4_io_in_a_Im = io_in_4_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_clock = clock;
  assign FPComplexMult_reducable_v2_5_reset = reset;
  assign FPComplexMult_reducable_v2_5_io_in_a_Re = io_in_5_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_io_in_a_Im = io_in_5_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_6_clock = clock;
  assign FPComplexMult_reducable_v2_6_reset = reset;
  assign FPComplexMult_reducable_v2_6_io_in_a_Re = io_in_6_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_6_io_in_a_Im = io_in_6_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_clock = clock;
  assign FPComplexMult_reducable_v2_7_reset = reset;
  assign FPComplexMult_reducable_v2_7_io_in_a_Re = io_in_7_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_io_in_a_Im = io_in_7_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_8_clock = clock;
  assign FPComplexMult_reducable_v2_8_reset = reset;
  assign FPComplexMult_reducable_v2_8_io_in_a_Re = io_in_8_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_8_io_in_a_Im = io_in_8_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_clock = clock;
  assign FPComplexMult_reducable_v2_9_reset = reset;
  assign FPComplexMult_reducable_v2_9_io_in_a_Re = io_in_9_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_io_in_a_Im = io_in_9_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_9_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_10_clock = clock;
  assign FPComplexMult_reducable_v2_10_reset = reset;
  assign FPComplexMult_reducable_v2_10_io_in_a_Re = io_in_10_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_10_io_in_a_Im = io_in_10_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_clock = clock;
  assign FPComplexMult_reducable_v2_11_reset = reset;
  assign FPComplexMult_reducable_v2_11_io_in_a_Re = io_in_11_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_io_in_a_Im = io_in_11_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_11_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_12_clock = clock;
  assign FPComplexMult_reducable_v2_12_reset = reset;
  assign FPComplexMult_reducable_v2_12_io_in_a_Re = io_in_12_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_12_io_in_a_Im = io_in_12_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_clock = clock;
  assign FPComplexMult_reducable_v2_13_reset = reset;
  assign FPComplexMult_reducable_v2_13_io_in_a_Re = io_in_13_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_io_in_a_Im = io_in_13_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_13_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_14_clock = clock;
  assign FPComplexMult_reducable_v2_14_reset = reset;
  assign FPComplexMult_reducable_v2_14_io_in_a_Re = io_in_14_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_14_io_in_a_Im = io_in_14_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_clock = clock;
  assign FPComplexMult_reducable_v2_15_reset = reset;
  assign FPComplexMult_reducable_v2_15_io_in_a_Re = io_in_15_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_io_in_a_Im = io_in_15_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_15_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_16_clock = clock;
  assign FPComplexMult_reducable_v2_16_reset = reset;
  assign FPComplexMult_reducable_v2_16_io_in_a_Re = io_in_16_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_16_io_in_a_Im = io_in_16_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_17_clock = clock;
  assign FPComplexMult_reducable_v2_17_reset = reset;
  assign FPComplexMult_reducable_v2_17_io_in_a_Re = io_in_17_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_17_io_in_a_Im = io_in_17_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_18_clock = clock;
  assign FPComplexMult_reducable_v2_18_reset = reset;
  assign FPComplexMult_reducable_v2_18_io_in_a_Re = io_in_18_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_18_io_in_a_Im = io_in_18_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_clock = clock;
  assign FPComplexMult_reducable_v2_19_reset = reset;
  assign FPComplexMult_reducable_v2_19_io_in_a_Re = io_in_19_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_io_in_a_Im = io_in_19_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_20_clock = clock;
  assign FPComplexMult_reducable_v2_20_reset = reset;
  assign FPComplexMult_reducable_v2_20_io_in_a_Re = io_in_20_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_20_io_in_a_Im = io_in_20_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_clock = clock;
  assign FPComplexMult_reducable_v2_21_reset = reset;
  assign FPComplexMult_reducable_v2_21_io_in_a_Re = io_in_21_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_io_in_a_Im = io_in_21_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_22_clock = clock;
  assign FPComplexMult_reducable_v2_22_reset = reset;
  assign FPComplexMult_reducable_v2_22_io_in_a_Re = io_in_22_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_22_io_in_a_Im = io_in_22_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_clock = clock;
  assign FPComplexMult_reducable_v2_23_reset = reset;
  assign FPComplexMult_reducable_v2_23_io_in_a_Re = io_in_23_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_io_in_a_Im = io_in_23_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_24_clock = clock;
  assign FPComplexMult_reducable_v2_24_reset = reset;
  assign FPComplexMult_reducable_v2_24_io_in_a_Re = io_in_24_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_24_io_in_a_Im = io_in_24_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_clock = clock;
  assign FPComplexMult_reducable_v2_25_reset = reset;
  assign FPComplexMult_reducable_v2_25_io_in_a_Re = io_in_25_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_io_in_a_Im = io_in_25_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_25_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_26_clock = clock;
  assign FPComplexMult_reducable_v2_26_reset = reset;
  assign FPComplexMult_reducable_v2_26_io_in_a_Re = io_in_26_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_26_io_in_a_Im = io_in_26_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_clock = clock;
  assign FPComplexMult_reducable_v2_27_reset = reset;
  assign FPComplexMult_reducable_v2_27_io_in_a_Re = io_in_27_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_io_in_a_Im = io_in_27_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_27_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_28_clock = clock;
  assign FPComplexMult_reducable_v2_28_reset = reset;
  assign FPComplexMult_reducable_v2_28_io_in_a_Re = io_in_28_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_28_io_in_a_Im = io_in_28_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_clock = clock;
  assign FPComplexMult_reducable_v2_29_reset = reset;
  assign FPComplexMult_reducable_v2_29_io_in_a_Re = io_in_29_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_io_in_a_Im = io_in_29_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_29_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_30_clock = clock;
  assign FPComplexMult_reducable_v2_30_reset = reset;
  assign FPComplexMult_reducable_v2_30_io_in_a_Re = io_in_30_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_30_io_in_a_Im = io_in_30_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_clock = clock;
  assign FPComplexMult_reducable_v2_31_reset = reset;
  assign FPComplexMult_reducable_v2_31_io_in_a_Re = io_in_31_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_io_in_a_Im = io_in_31_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_31_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
endmodule
module TwiddleFactors_2(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im
);
  wire  FPComplexMult_reducable_v2_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_1_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_1_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_2_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_2_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_3_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_3_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_4_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_4_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_5_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_5_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_6_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_6_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_7_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_7_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_8_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_8_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_9_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_9_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_10_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_10_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_11_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_11_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_12_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_12_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_13_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_13_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_14_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_14_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_15_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_15_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_16_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_16_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_17_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_17_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_18_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_18_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_19_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_19_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_20_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_20_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_21_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_21_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_22_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_22_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_23_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_23_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_24_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_24_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_25_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_25_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_26_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_26_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_27_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_27_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_28_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_28_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_29_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_29_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_30_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_30_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_31_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_31_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_clock),
    .reset(FPComplexMult_reducable_v2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_1 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_1_clock),
    .reset(FPComplexMult_reducable_v2_1_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_1_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_1_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_2 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_2_clock),
    .reset(FPComplexMult_reducable_v2_2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_3 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_3_clock),
    .reset(FPComplexMult_reducable_v2_3_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_3_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_3_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_4 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_4_clock),
    .reset(FPComplexMult_reducable_v2_4_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_4_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_4_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_5 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_5_clock),
    .reset(FPComplexMult_reducable_v2_5_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_5_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_6 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_6_clock),
    .reset(FPComplexMult_reducable_v2_6_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_6_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_6_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_7 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_7_clock),
    .reset(FPComplexMult_reducable_v2_7_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_7_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_8 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_8_clock),
    .reset(FPComplexMult_reducable_v2_8_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_8_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_8_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_9 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_9_clock),
    .reset(FPComplexMult_reducable_v2_9_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_9_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_10 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_10_clock),
    .reset(FPComplexMult_reducable_v2_10_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_10_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_10_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_11 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_11_clock),
    .reset(FPComplexMult_reducable_v2_11_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_11_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_12 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_12_clock),
    .reset(FPComplexMult_reducable_v2_12_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_12_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_12_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_13 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_13_clock),
    .reset(FPComplexMult_reducable_v2_13_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_13_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_14 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_14_clock),
    .reset(FPComplexMult_reducable_v2_14_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_14_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_14_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_15 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_15_clock),
    .reset(FPComplexMult_reducable_v2_15_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_15_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_16 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_16_clock),
    .reset(FPComplexMult_reducable_v2_16_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_16_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_16_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_16_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_16_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_113 FPComplexMult_reducable_v2_17 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_17_clock),
    .reset(FPComplexMult_reducable_v2_17_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_17_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_17_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_17_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_17_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_18 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_18_clock),
    .reset(FPComplexMult_reducable_v2_18_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_18_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_18_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_18_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_18_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_113 FPComplexMult_reducable_v2_19 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_19_clock),
    .reset(FPComplexMult_reducable_v2_19_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_19_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_19_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_19_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_19_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_20 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_20_clock),
    .reset(FPComplexMult_reducable_v2_20_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_20_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_20_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_20_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_20_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_21 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_21_clock),
    .reset(FPComplexMult_reducable_v2_21_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_21_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_21_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_21_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_21_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_21_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_21_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_22 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_22_clock),
    .reset(FPComplexMult_reducable_v2_22_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_22_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_22_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_22_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_22_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_23 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_23_clock),
    .reset(FPComplexMult_reducable_v2_23_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_23_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_23_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_23_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_23_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_23_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_23_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_24 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_24_clock),
    .reset(FPComplexMult_reducable_v2_24_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_24_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_24_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_24_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_24_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_25 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_25_clock),
    .reset(FPComplexMult_reducable_v2_25_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_25_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_25_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_25_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_25_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_25_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_25_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_26 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_26_clock),
    .reset(FPComplexMult_reducable_v2_26_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_26_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_26_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_26_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_26_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_27 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_27_clock),
    .reset(FPComplexMult_reducable_v2_27_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_27_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_27_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_27_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_27_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_27_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_27_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_28 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_28_clock),
    .reset(FPComplexMult_reducable_v2_28_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_28_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_28_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_28_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_28_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_29 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_29_clock),
    .reset(FPComplexMult_reducable_v2_29_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_29_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_29_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_29_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_29_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_29_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_29_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_30 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_30_clock),
    .reset(FPComplexMult_reducable_v2_30_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_30_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_30_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_30_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_30_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_31 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_31_clock),
    .reset(FPComplexMult_reducable_v2_31_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_31_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_31_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_31_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_31_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_31_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_31_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_0_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_1_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_1_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_2_Re = FPComplexMult_reducable_v2_2_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_2_Im = FPComplexMult_reducable_v2_2_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_3_Re = FPComplexMult_reducable_v2_3_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_3_Im = FPComplexMult_reducable_v2_3_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_4_Re = FPComplexMult_reducable_v2_4_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_4_Im = FPComplexMult_reducable_v2_4_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_5_Re = FPComplexMult_reducable_v2_5_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_5_Im = FPComplexMult_reducable_v2_5_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_6_Re = FPComplexMult_reducable_v2_6_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_6_Im = FPComplexMult_reducable_v2_6_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_7_Re = FPComplexMult_reducable_v2_7_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_7_Im = FPComplexMult_reducable_v2_7_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_8_Re = FPComplexMult_reducable_v2_8_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_8_Im = FPComplexMult_reducable_v2_8_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_9_Re = FPComplexMult_reducable_v2_9_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_9_Im = FPComplexMult_reducable_v2_9_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_10_Re = FPComplexMult_reducable_v2_10_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_10_Im = FPComplexMult_reducable_v2_10_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_11_Re = FPComplexMult_reducable_v2_11_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_11_Im = FPComplexMult_reducable_v2_11_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_12_Re = FPComplexMult_reducable_v2_12_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_12_Im = FPComplexMult_reducable_v2_12_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_13_Re = FPComplexMult_reducable_v2_13_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_13_Im = FPComplexMult_reducable_v2_13_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_14_Re = FPComplexMult_reducable_v2_14_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_14_Im = FPComplexMult_reducable_v2_14_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_15_Re = FPComplexMult_reducable_v2_15_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_15_Im = FPComplexMult_reducable_v2_15_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_16_Re = FPComplexMult_reducable_v2_16_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_16_Im = FPComplexMult_reducable_v2_16_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_17_Re = FPComplexMult_reducable_v2_17_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_17_Im = FPComplexMult_reducable_v2_17_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_18_Re = FPComplexMult_reducable_v2_18_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_18_Im = FPComplexMult_reducable_v2_18_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_19_Re = FPComplexMult_reducable_v2_19_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_19_Im = FPComplexMult_reducable_v2_19_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_20_Re = FPComplexMult_reducable_v2_20_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_20_Im = FPComplexMult_reducable_v2_20_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_21_Re = FPComplexMult_reducable_v2_21_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_21_Im = FPComplexMult_reducable_v2_21_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_22_Re = FPComplexMult_reducable_v2_22_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_22_Im = FPComplexMult_reducable_v2_22_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_23_Re = FPComplexMult_reducable_v2_23_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_23_Im = FPComplexMult_reducable_v2_23_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_24_Re = FPComplexMult_reducable_v2_24_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_24_Im = FPComplexMult_reducable_v2_24_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_25_Re = FPComplexMult_reducable_v2_25_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_25_Im = FPComplexMult_reducable_v2_25_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_26_Re = FPComplexMult_reducable_v2_26_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_26_Im = FPComplexMult_reducable_v2_26_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_27_Re = FPComplexMult_reducable_v2_27_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_27_Im = FPComplexMult_reducable_v2_27_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_28_Re = FPComplexMult_reducable_v2_28_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_28_Im = FPComplexMult_reducable_v2_28_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_29_Re = FPComplexMult_reducable_v2_29_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_29_Im = FPComplexMult_reducable_v2_29_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_30_Re = FPComplexMult_reducable_v2_30_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_30_Im = FPComplexMult_reducable_v2_30_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_31_Re = FPComplexMult_reducable_v2_31_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_31_Im = FPComplexMult_reducable_v2_31_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign FPComplexMult_reducable_v2_clock = clock;
  assign FPComplexMult_reducable_v2_reset = reset;
  assign FPComplexMult_reducable_v2_io_in_a_Re = io_in_0_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_io_in_a_Im = io_in_0_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_1_clock = clock;
  assign FPComplexMult_reducable_v2_1_reset = reset;
  assign FPComplexMult_reducable_v2_1_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_1_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_2_clock = clock;
  assign FPComplexMult_reducable_v2_2_reset = reset;
  assign FPComplexMult_reducable_v2_2_io_in_a_Re = io_in_2_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_2_io_in_a_Im = io_in_2_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_clock = clock;
  assign FPComplexMult_reducable_v2_3_reset = reset;
  assign FPComplexMult_reducable_v2_3_io_in_a_Re = io_in_3_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_io_in_a_Im = io_in_3_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_4_clock = clock;
  assign FPComplexMult_reducable_v2_4_reset = reset;
  assign FPComplexMult_reducable_v2_4_io_in_a_Re = io_in_4_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_4_io_in_a_Im = io_in_4_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_clock = clock;
  assign FPComplexMult_reducable_v2_5_reset = reset;
  assign FPComplexMult_reducable_v2_5_io_in_a_Re = io_in_5_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_io_in_a_Im = io_in_5_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_io_in_b_Re = 32'h3f6c835e; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_5_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_6_clock = clock;
  assign FPComplexMult_reducable_v2_6_reset = reset;
  assign FPComplexMult_reducable_v2_6_io_in_a_Re = io_in_6_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_6_io_in_a_Im = io_in_6_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_clock = clock;
  assign FPComplexMult_reducable_v2_7_reset = reset;
  assign FPComplexMult_reducable_v2_7_io_in_a_Re = io_in_7_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_io_in_a_Im = io_in_7_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_io_in_b_Re = 32'h3f6c835e; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_7_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_8_clock = clock;
  assign FPComplexMult_reducable_v2_8_reset = reset;
  assign FPComplexMult_reducable_v2_8_io_in_a_Re = io_in_8_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_8_io_in_a_Im = io_in_8_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_clock = clock;
  assign FPComplexMult_reducable_v2_9_reset = reset;
  assign FPComplexMult_reducable_v2_9_io_in_a_Re = io_in_9_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_io_in_a_Im = io_in_9_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_9_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_10_clock = clock;
  assign FPComplexMult_reducable_v2_10_reset = reset;
  assign FPComplexMult_reducable_v2_10_io_in_a_Re = io_in_10_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_10_io_in_a_Im = io_in_10_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_clock = clock;
  assign FPComplexMult_reducable_v2_11_reset = reset;
  assign FPComplexMult_reducable_v2_11_io_in_a_Re = io_in_11_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_io_in_a_Im = io_in_11_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_11_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_12_clock = clock;
  assign FPComplexMult_reducable_v2_12_reset = reset;
  assign FPComplexMult_reducable_v2_12_io_in_a_Re = io_in_12_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_12_io_in_a_Im = io_in_12_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_clock = clock;
  assign FPComplexMult_reducable_v2_13_reset = reset;
  assign FPComplexMult_reducable_v2_13_io_in_a_Re = io_in_13_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_io_in_a_Im = io_in_13_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_io_in_b_Re = 32'h3ec3ef14; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_13_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_14_clock = clock;
  assign FPComplexMult_reducable_v2_14_reset = reset;
  assign FPComplexMult_reducable_v2_14_io_in_a_Re = io_in_14_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_14_io_in_a_Im = io_in_14_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_clock = clock;
  assign FPComplexMult_reducable_v2_15_reset = reset;
  assign FPComplexMult_reducable_v2_15_io_in_a_Re = io_in_15_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_io_in_a_Im = io_in_15_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_io_in_b_Re = 32'h3ec3ef14; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_15_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_16_clock = clock;
  assign FPComplexMult_reducable_v2_16_reset = reset;
  assign FPComplexMult_reducable_v2_16_io_in_a_Re = io_in_16_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_16_io_in_a_Im = io_in_16_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_17_clock = clock;
  assign FPComplexMult_reducable_v2_17_reset = reset;
  assign FPComplexMult_reducable_v2_17_io_in_a_Re = io_in_17_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_17_io_in_a_Im = io_in_17_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_18_clock = clock;
  assign FPComplexMult_reducable_v2_18_reset = reset;
  assign FPComplexMult_reducable_v2_18_io_in_a_Re = io_in_18_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_18_io_in_a_Im = io_in_18_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_clock = clock;
  assign FPComplexMult_reducable_v2_19_reset = reset;
  assign FPComplexMult_reducable_v2_19_io_in_a_Re = io_in_19_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_io_in_a_Im = io_in_19_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_20_clock = clock;
  assign FPComplexMult_reducable_v2_20_reset = reset;
  assign FPComplexMult_reducable_v2_20_io_in_a_Re = io_in_20_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_20_io_in_a_Im = io_in_20_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_clock = clock;
  assign FPComplexMult_reducable_v2_21_reset = reset;
  assign FPComplexMult_reducable_v2_21_io_in_a_Re = io_in_21_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_io_in_a_Im = io_in_21_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_io_in_b_Re = 32'hbec3ef14; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_21_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_22_clock = clock;
  assign FPComplexMult_reducable_v2_22_reset = reset;
  assign FPComplexMult_reducable_v2_22_io_in_a_Re = io_in_22_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_22_io_in_a_Im = io_in_22_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_clock = clock;
  assign FPComplexMult_reducable_v2_23_reset = reset;
  assign FPComplexMult_reducable_v2_23_io_in_a_Re = io_in_23_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_io_in_a_Im = io_in_23_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_io_in_b_Re = 32'hbec3ef14; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_23_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_24_clock = clock;
  assign FPComplexMult_reducable_v2_24_reset = reset;
  assign FPComplexMult_reducable_v2_24_io_in_a_Re = io_in_24_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_24_io_in_a_Im = io_in_24_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_clock = clock;
  assign FPComplexMult_reducable_v2_25_reset = reset;
  assign FPComplexMult_reducable_v2_25_io_in_a_Re = io_in_25_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_io_in_a_Im = io_in_25_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_25_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_26_clock = clock;
  assign FPComplexMult_reducable_v2_26_reset = reset;
  assign FPComplexMult_reducable_v2_26_io_in_a_Re = io_in_26_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_26_io_in_a_Im = io_in_26_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_clock = clock;
  assign FPComplexMult_reducable_v2_27_reset = reset;
  assign FPComplexMult_reducable_v2_27_io_in_a_Re = io_in_27_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_io_in_a_Im = io_in_27_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_27_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_28_clock = clock;
  assign FPComplexMult_reducable_v2_28_reset = reset;
  assign FPComplexMult_reducable_v2_28_io_in_a_Re = io_in_28_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_28_io_in_a_Im = io_in_28_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_clock = clock;
  assign FPComplexMult_reducable_v2_29_reset = reset;
  assign FPComplexMult_reducable_v2_29_io_in_a_Re = io_in_29_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_io_in_a_Im = io_in_29_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_io_in_b_Re = 32'hbf6c835e; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_29_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_30_clock = clock;
  assign FPComplexMult_reducable_v2_30_reset = reset;
  assign FPComplexMult_reducable_v2_30_io_in_a_Re = io_in_30_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_30_io_in_a_Im = io_in_30_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_clock = clock;
  assign FPComplexMult_reducable_v2_31_reset = reset;
  assign FPComplexMult_reducable_v2_31_io_in_a_Re = io_in_31_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_io_in_a_Im = io_in_31_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_io_in_b_Re = 32'hbf6c835e; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_31_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 2304:30]
endmodule
module TwiddleFactors_3(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im
);
  wire  FPComplexMult_reducable_v2_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_1_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_1_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_2_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_2_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_2_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_3_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_3_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_3_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_4_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_4_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_4_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_5_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_5_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_5_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_6_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_6_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_6_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_7_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_7_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_7_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_8_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_8_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_8_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_9_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_9_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_9_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_10_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_10_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_10_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_11_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_11_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_11_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_12_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_12_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_12_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_13_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_13_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_13_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_14_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_14_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_14_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_15_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_15_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_15_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_16_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_16_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_16_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_17_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_17_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_17_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_18_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_18_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_18_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_19_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_19_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_19_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_20_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_20_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_20_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_21_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_21_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_21_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_22_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_22_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_22_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_23_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_23_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_23_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_24_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_24_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_24_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_25_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_25_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_25_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_26_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_26_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_26_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_27_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_27_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_27_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_28_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_28_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_28_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_29_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_29_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_29_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_30_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_30_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_30_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_31_clock; // @[FFTDesigns.scala 2298:28]
  wire  FPComplexMult_reducable_v2_31_reset; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_a_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_a_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_b_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_in_b_Im; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_out_s_Re; // @[FFTDesigns.scala 2298:28]
  wire [31:0] FPComplexMult_reducable_v2_31_io_out_s_Im; // @[FFTDesigns.scala 2298:28]
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_clock),
    .reset(FPComplexMult_reducable_v2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_1 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_1_clock),
    .reset(FPComplexMult_reducable_v2_1_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_1_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_1_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_2 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_2_clock),
    .reset(FPComplexMult_reducable_v2_2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_3 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_3_clock),
    .reset(FPComplexMult_reducable_v2_3_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_3_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_4 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_4_clock),
    .reset(FPComplexMult_reducable_v2_4_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_4_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_4_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_5 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_5_clock),
    .reset(FPComplexMult_reducable_v2_5_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_5_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_6 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_6_clock),
    .reset(FPComplexMult_reducable_v2_6_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_6_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_6_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_7 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_7_clock),
    .reset(FPComplexMult_reducable_v2_7_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_7_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_8 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_8_clock),
    .reset(FPComplexMult_reducable_v2_8_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_8_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_8_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_9 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_9_clock),
    .reset(FPComplexMult_reducable_v2_9_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_9_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_10 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_10_clock),
    .reset(FPComplexMult_reducable_v2_10_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_10_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_10_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_11 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_11_clock),
    .reset(FPComplexMult_reducable_v2_11_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_11_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_12 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_12_clock),
    .reset(FPComplexMult_reducable_v2_12_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_12_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_12_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_13 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_13_clock),
    .reset(FPComplexMult_reducable_v2_13_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_13_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_14 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_14_clock),
    .reset(FPComplexMult_reducable_v2_14_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_14_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_14_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_15 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_15_clock),
    .reset(FPComplexMult_reducable_v2_15_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_15_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_16 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_16_clock),
    .reset(FPComplexMult_reducable_v2_16_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_16_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_16_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_16_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_16_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_113 FPComplexMult_reducable_v2_17 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_17_clock),
    .reset(FPComplexMult_reducable_v2_17_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_17_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_17_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_17_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_17_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_18 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_18_clock),
    .reset(FPComplexMult_reducable_v2_18_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_18_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_18_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_18_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_18_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_19 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_19_clock),
    .reset(FPComplexMult_reducable_v2_19_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_19_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_19_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_19_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_19_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_19_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_19_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_20 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_20_clock),
    .reset(FPComplexMult_reducable_v2_20_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_20_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_20_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_20_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_20_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_21 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_21_clock),
    .reset(FPComplexMult_reducable_v2_21_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_21_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_21_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_21_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_21_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_21_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_21_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_22 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_22_clock),
    .reset(FPComplexMult_reducable_v2_22_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_22_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_22_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_22_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_22_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_23 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_23_clock),
    .reset(FPComplexMult_reducable_v2_23_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_23_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_23_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_23_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_23_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_23_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_23_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_24 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_24_clock),
    .reset(FPComplexMult_reducable_v2_24_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_24_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_24_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_24_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_24_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_25 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_25_clock),
    .reset(FPComplexMult_reducable_v2_25_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_25_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_25_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_25_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_25_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_25_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_25_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_26 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_26_clock),
    .reset(FPComplexMult_reducable_v2_26_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_26_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_26_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_26_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_26_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_27 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_27_clock),
    .reset(FPComplexMult_reducable_v2_27_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_27_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_27_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_27_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_27_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_27_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_27_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_28 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_28_clock),
    .reset(FPComplexMult_reducable_v2_28_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_28_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_28_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_28_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_28_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_29 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_29_clock),
    .reset(FPComplexMult_reducable_v2_29_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_29_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_29_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_29_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_29_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_29_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_29_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_96 FPComplexMult_reducable_v2_30 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_30_clock),
    .reset(FPComplexMult_reducable_v2_30_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_30_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_30_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_30_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_30_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_v2_31 ( // @[FFTDesigns.scala 2298:28]
    .clock(FPComplexMult_reducable_v2_31_clock),
    .reset(FPComplexMult_reducable_v2_31_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_31_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_31_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_v2_31_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_v2_31_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_31_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_31_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_0_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_1_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_1_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_2_Re = FPComplexMult_reducable_v2_2_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_2_Im = FPComplexMult_reducable_v2_2_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_3_Re = FPComplexMult_reducable_v2_3_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_3_Im = FPComplexMult_reducable_v2_3_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_4_Re = FPComplexMult_reducable_v2_4_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_4_Im = FPComplexMult_reducable_v2_4_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_5_Re = FPComplexMult_reducable_v2_5_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_5_Im = FPComplexMult_reducable_v2_5_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_6_Re = FPComplexMult_reducable_v2_6_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_6_Im = FPComplexMult_reducable_v2_6_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_7_Re = FPComplexMult_reducable_v2_7_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_7_Im = FPComplexMult_reducable_v2_7_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_8_Re = FPComplexMult_reducable_v2_8_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_8_Im = FPComplexMult_reducable_v2_8_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_9_Re = FPComplexMult_reducable_v2_9_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_9_Im = FPComplexMult_reducable_v2_9_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_10_Re = FPComplexMult_reducable_v2_10_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_10_Im = FPComplexMult_reducable_v2_10_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_11_Re = FPComplexMult_reducable_v2_11_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_11_Im = FPComplexMult_reducable_v2_11_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_12_Re = FPComplexMult_reducable_v2_12_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_12_Im = FPComplexMult_reducable_v2_12_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_13_Re = FPComplexMult_reducable_v2_13_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_13_Im = FPComplexMult_reducable_v2_13_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_14_Re = FPComplexMult_reducable_v2_14_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_14_Im = FPComplexMult_reducable_v2_14_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_15_Re = FPComplexMult_reducable_v2_15_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_15_Im = FPComplexMult_reducable_v2_15_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_16_Re = FPComplexMult_reducable_v2_16_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_16_Im = FPComplexMult_reducable_v2_16_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_17_Re = FPComplexMult_reducable_v2_17_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_17_Im = FPComplexMult_reducable_v2_17_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_18_Re = FPComplexMult_reducable_v2_18_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_18_Im = FPComplexMult_reducable_v2_18_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_19_Re = FPComplexMult_reducable_v2_19_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_19_Im = FPComplexMult_reducable_v2_19_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_20_Re = FPComplexMult_reducable_v2_20_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_20_Im = FPComplexMult_reducable_v2_20_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_21_Re = FPComplexMult_reducable_v2_21_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_21_Im = FPComplexMult_reducable_v2_21_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_22_Re = FPComplexMult_reducable_v2_22_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_22_Im = FPComplexMult_reducable_v2_22_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_23_Re = FPComplexMult_reducable_v2_23_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_23_Im = FPComplexMult_reducable_v2_23_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_24_Re = FPComplexMult_reducable_v2_24_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_24_Im = FPComplexMult_reducable_v2_24_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_25_Re = FPComplexMult_reducable_v2_25_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_25_Im = FPComplexMult_reducable_v2_25_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_26_Re = FPComplexMult_reducable_v2_26_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_26_Im = FPComplexMult_reducable_v2_26_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_27_Re = FPComplexMult_reducable_v2_27_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_27_Im = FPComplexMult_reducable_v2_27_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_28_Re = FPComplexMult_reducable_v2_28_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_28_Im = FPComplexMult_reducable_v2_28_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_29_Re = FPComplexMult_reducable_v2_29_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_29_Im = FPComplexMult_reducable_v2_29_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_30_Re = FPComplexMult_reducable_v2_30_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_30_Im = FPComplexMult_reducable_v2_30_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign io_out_31_Re = FPComplexMult_reducable_v2_31_io_out_s_Re; // @[FFTDesigns.scala 2305:17]
  assign io_out_31_Im = FPComplexMult_reducable_v2_31_io_out_s_Im; // @[FFTDesigns.scala 2305:17]
  assign FPComplexMult_reducable_v2_clock = clock;
  assign FPComplexMult_reducable_v2_reset = reset;
  assign FPComplexMult_reducable_v2_io_in_a_Re = io_in_0_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_io_in_a_Im = io_in_0_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_1_clock = clock;
  assign FPComplexMult_reducable_v2_1_reset = reset;
  assign FPComplexMult_reducable_v2_1_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_1_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_2_clock = clock;
  assign FPComplexMult_reducable_v2_2_reset = reset;
  assign FPComplexMult_reducable_v2_2_io_in_a_Re = io_in_2_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_2_io_in_a_Im = io_in_2_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_clock = clock;
  assign FPComplexMult_reducable_v2_3_reset = reset;
  assign FPComplexMult_reducable_v2_3_io_in_a_Re = io_in_3_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_io_in_a_Im = io_in_3_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_3_io_in_b_Re = 32'h3f7b14be; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_3_io_in_b_Im = 32'hbe47c5c0; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_4_clock = clock;
  assign FPComplexMult_reducable_v2_4_reset = reset;
  assign FPComplexMult_reducable_v2_4_io_in_a_Re = io_in_4_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_4_io_in_a_Im = io_in_4_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_clock = clock;
  assign FPComplexMult_reducable_v2_5_reset = reset;
  assign FPComplexMult_reducable_v2_5_io_in_a_Re = io_in_5_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_io_in_a_Im = io_in_5_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_5_io_in_b_Re = 32'h3f6c835e; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_5_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_6_clock = clock;
  assign FPComplexMult_reducable_v2_6_reset = reset;
  assign FPComplexMult_reducable_v2_6_io_in_a_Re = io_in_6_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_6_io_in_a_Im = io_in_6_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_clock = clock;
  assign FPComplexMult_reducable_v2_7_reset = reset;
  assign FPComplexMult_reducable_v2_7_io_in_a_Re = io_in_7_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_io_in_a_Im = io_in_7_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_7_io_in_b_Re = 32'h3f54db30; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_7_io_in_b_Im = 32'hbf0e39d8; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_8_clock = clock;
  assign FPComplexMult_reducable_v2_8_reset = reset;
  assign FPComplexMult_reducable_v2_8_io_in_a_Re = io_in_8_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_8_io_in_a_Im = io_in_8_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_clock = clock;
  assign FPComplexMult_reducable_v2_9_reset = reset;
  assign FPComplexMult_reducable_v2_9_io_in_a_Re = io_in_9_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_io_in_a_Im = io_in_9_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_9_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_9_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_10_clock = clock;
  assign FPComplexMult_reducable_v2_10_reset = reset;
  assign FPComplexMult_reducable_v2_10_io_in_a_Re = io_in_10_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_10_io_in_a_Im = io_in_10_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_clock = clock;
  assign FPComplexMult_reducable_v2_11_reset = reset;
  assign FPComplexMult_reducable_v2_11_io_in_a_Re = io_in_11_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_io_in_a_Im = io_in_11_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_11_io_in_b_Re = 32'h3f0e39d8; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_11_io_in_b_Im = 32'hbf54db30; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_12_clock = clock;
  assign FPComplexMult_reducable_v2_12_reset = reset;
  assign FPComplexMult_reducable_v2_12_io_in_a_Re = io_in_12_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_12_io_in_a_Im = io_in_12_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_clock = clock;
  assign FPComplexMult_reducable_v2_13_reset = reset;
  assign FPComplexMult_reducable_v2_13_io_in_a_Re = io_in_13_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_io_in_a_Im = io_in_13_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_13_io_in_b_Re = 32'h3ec3ef14; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_13_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_14_clock = clock;
  assign FPComplexMult_reducable_v2_14_reset = reset;
  assign FPComplexMult_reducable_v2_14_io_in_a_Re = io_in_14_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_14_io_in_a_Im = io_in_14_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_clock = clock;
  assign FPComplexMult_reducable_v2_15_reset = reset;
  assign FPComplexMult_reducable_v2_15_io_in_a_Re = io_in_15_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_io_in_a_Im = io_in_15_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_15_io_in_b_Re = 32'h3e47c5c0; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_15_io_in_b_Im = 32'hbf7b14be; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_16_clock = clock;
  assign FPComplexMult_reducable_v2_16_reset = reset;
  assign FPComplexMult_reducable_v2_16_io_in_a_Re = io_in_16_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_16_io_in_a_Im = io_in_16_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_17_clock = clock;
  assign FPComplexMult_reducable_v2_17_reset = reset;
  assign FPComplexMult_reducable_v2_17_io_in_a_Re = io_in_17_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_17_io_in_a_Im = io_in_17_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_18_clock = clock;
  assign FPComplexMult_reducable_v2_18_reset = reset;
  assign FPComplexMult_reducable_v2_18_io_in_a_Re = io_in_18_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_18_io_in_a_Im = io_in_18_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_clock = clock;
  assign FPComplexMult_reducable_v2_19_reset = reset;
  assign FPComplexMult_reducable_v2_19_io_in_a_Re = io_in_19_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_io_in_a_Im = io_in_19_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_19_io_in_b_Re = 32'hbe47c5c0; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_19_io_in_b_Im = 32'hbf7b14be; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_20_clock = clock;
  assign FPComplexMult_reducable_v2_20_reset = reset;
  assign FPComplexMult_reducable_v2_20_io_in_a_Re = io_in_20_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_20_io_in_a_Im = io_in_20_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_clock = clock;
  assign FPComplexMult_reducable_v2_21_reset = reset;
  assign FPComplexMult_reducable_v2_21_io_in_a_Re = io_in_21_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_io_in_a_Im = io_in_21_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_21_io_in_b_Re = 32'hbec3ef14; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_21_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_22_clock = clock;
  assign FPComplexMult_reducable_v2_22_reset = reset;
  assign FPComplexMult_reducable_v2_22_io_in_a_Re = io_in_22_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_22_io_in_a_Im = io_in_22_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_clock = clock;
  assign FPComplexMult_reducable_v2_23_reset = reset;
  assign FPComplexMult_reducable_v2_23_io_in_a_Re = io_in_23_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_io_in_a_Im = io_in_23_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_23_io_in_b_Re = 32'hbf0e39d8; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_23_io_in_b_Im = 32'hbf54db30; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_24_clock = clock;
  assign FPComplexMult_reducable_v2_24_reset = reset;
  assign FPComplexMult_reducable_v2_24_io_in_a_Re = io_in_24_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_24_io_in_a_Im = io_in_24_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_clock = clock;
  assign FPComplexMult_reducable_v2_25_reset = reset;
  assign FPComplexMult_reducable_v2_25_io_in_a_Re = io_in_25_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_io_in_a_Im = io_in_25_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_25_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_25_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_26_clock = clock;
  assign FPComplexMult_reducable_v2_26_reset = reset;
  assign FPComplexMult_reducable_v2_26_io_in_a_Re = io_in_26_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_26_io_in_a_Im = io_in_26_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_clock = clock;
  assign FPComplexMult_reducable_v2_27_reset = reset;
  assign FPComplexMult_reducable_v2_27_io_in_a_Re = io_in_27_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_io_in_a_Im = io_in_27_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_27_io_in_b_Re = 32'hbf54db30; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_27_io_in_b_Im = 32'hbf0e39d8; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_28_clock = clock;
  assign FPComplexMult_reducable_v2_28_reset = reset;
  assign FPComplexMult_reducable_v2_28_io_in_a_Re = io_in_28_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_28_io_in_a_Im = io_in_28_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_clock = clock;
  assign FPComplexMult_reducable_v2_29_reset = reset;
  assign FPComplexMult_reducable_v2_29_io_in_a_Re = io_in_29_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_io_in_a_Im = io_in_29_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_29_io_in_b_Re = 32'hbf6c835e; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_29_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 2304:30]
  assign FPComplexMult_reducable_v2_30_clock = clock;
  assign FPComplexMult_reducable_v2_30_reset = reset;
  assign FPComplexMult_reducable_v2_30_io_in_a_Re = io_in_30_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_30_io_in_a_Im = io_in_30_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_clock = clock;
  assign FPComplexMult_reducable_v2_31_reset = reset;
  assign FPComplexMult_reducable_v2_31_io_in_a_Re = io_in_31_Re; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_io_in_a_Im = io_in_31_Im; // @[FFTDesigns.scala 2302:27]
  assign FPComplexMult_reducable_v2_31_io_in_b_Re = 32'hbf7b14be; // @[FFTDesigns.scala 2303:30]
  assign FPComplexMult_reducable_v2_31_io_in_b_Im = 32'hbe47c5c0; // @[FFTDesigns.scala 2304:30]
endmodule
module FFT_sr_v2_nrv_32(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im
);
  wire  DFT_r_v2_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_1_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_1_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_1_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_1_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_1_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_1_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_2_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_2_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_2_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_2_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_2_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_2_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_3_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_3_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_3_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_3_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_3_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_3_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_4_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_4_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_4_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_4_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_4_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_4_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_4_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_4_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_4_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_4_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_5_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_5_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_5_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_5_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_5_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_5_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_5_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_5_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_5_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_5_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_6_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_6_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_6_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_6_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_6_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_6_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_6_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_6_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_6_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_6_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_7_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_7_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_7_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_7_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_7_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_7_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_7_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_7_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_7_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_7_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_8_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_8_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_8_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_8_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_8_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_8_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_8_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_8_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_8_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_8_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_9_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_9_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_9_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_9_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_9_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_9_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_9_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_9_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_9_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_9_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_10_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_10_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_10_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_10_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_10_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_10_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_10_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_10_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_10_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_10_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_11_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_11_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_11_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_11_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_11_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_11_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_11_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_11_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_11_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_11_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_12_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_12_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_12_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_12_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_12_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_12_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_12_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_12_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_12_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_12_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_13_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_13_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_13_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_13_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_13_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_13_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_13_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_13_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_13_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_13_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_14_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_14_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_14_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_14_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_14_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_14_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_14_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_14_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_14_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_14_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_15_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_15_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_15_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_15_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_15_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_15_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_15_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_15_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_15_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_15_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_16_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_16_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_16_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_16_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_16_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_16_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_16_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_16_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_16_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_16_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_17_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_17_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_17_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_17_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_17_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_17_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_17_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_17_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_17_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_17_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_18_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_18_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_18_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_18_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_18_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_18_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_18_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_18_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_18_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_18_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_19_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_19_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_19_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_19_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_19_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_19_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_19_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_19_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_19_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_19_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_20_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_20_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_20_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_20_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_20_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_20_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_20_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_20_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_20_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_20_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_21_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_21_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_21_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_21_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_21_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_21_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_21_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_21_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_21_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_21_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_22_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_22_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_22_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_22_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_22_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_22_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_22_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_22_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_22_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_22_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_23_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_23_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_23_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_23_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_23_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_23_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_23_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_23_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_23_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_23_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_24_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_24_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_24_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_24_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_24_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_24_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_24_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_24_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_24_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_24_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_25_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_25_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_25_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_25_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_25_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_25_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_25_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_25_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_25_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_25_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_26_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_26_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_26_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_26_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_26_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_26_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_26_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_26_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_26_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_26_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_27_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_27_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_27_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_27_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_27_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_27_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_27_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_27_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_27_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_27_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_28_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_28_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_28_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_28_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_28_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_28_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_28_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_28_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_28_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_28_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_29_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_29_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_29_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_29_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_29_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_29_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_29_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_29_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_29_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_29_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_30_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_30_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_30_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_30_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_30_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_30_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_30_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_30_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_30_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_30_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_31_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_31_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_31_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_31_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_31_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_31_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_31_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_31_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_31_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_31_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_32_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_32_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_32_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_32_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_32_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_32_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_32_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_32_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_32_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_32_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_33_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_33_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_33_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_33_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_33_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_33_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_33_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_33_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_33_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_33_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_34_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_34_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_34_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_34_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_34_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_34_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_34_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_34_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_34_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_34_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_35_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_35_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_35_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_35_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_35_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_35_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_35_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_35_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_35_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_35_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_36_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_36_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_36_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_36_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_36_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_36_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_36_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_36_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_36_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_36_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_37_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_37_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_37_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_37_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_37_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_37_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_37_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_37_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_37_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_37_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_38_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_38_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_38_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_38_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_38_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_38_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_38_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_38_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_38_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_38_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_39_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_39_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_39_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_39_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_39_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_39_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_39_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_39_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_39_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_39_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_40_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_40_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_40_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_40_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_40_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_40_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_40_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_40_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_40_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_40_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_41_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_41_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_41_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_41_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_41_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_41_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_41_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_41_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_41_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_41_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_42_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_42_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_42_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_42_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_42_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_42_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_42_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_42_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_42_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_42_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_43_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_43_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_43_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_43_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_43_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_43_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_43_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_43_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_43_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_43_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_44_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_44_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_44_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_44_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_44_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_44_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_44_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_44_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_44_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_44_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_45_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_45_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_45_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_45_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_45_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_45_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_45_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_45_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_45_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_45_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_46_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_46_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_46_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_46_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_46_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_46_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_46_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_46_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_46_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_46_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_47_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_47_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_47_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_47_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_47_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_47_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_47_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_47_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_47_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_47_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_48_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_48_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_48_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_48_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_48_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_48_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_48_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_48_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_48_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_48_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_49_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_49_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_49_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_49_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_49_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_49_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_49_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_49_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_49_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_49_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_50_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_50_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_50_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_50_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_50_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_50_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_50_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_50_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_50_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_50_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_51_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_51_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_51_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_51_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_51_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_51_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_51_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_51_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_51_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_51_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_52_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_52_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_52_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_52_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_52_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_52_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_52_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_52_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_52_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_52_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_53_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_53_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_53_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_53_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_53_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_53_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_53_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_53_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_53_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_53_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_54_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_54_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_54_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_54_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_54_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_54_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_54_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_54_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_54_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_54_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_55_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_55_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_55_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_55_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_55_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_55_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_55_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_55_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_55_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_55_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_56_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_56_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_56_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_56_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_56_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_56_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_56_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_56_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_56_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_56_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_57_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_57_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_57_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_57_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_57_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_57_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_57_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_57_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_57_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_57_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_58_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_58_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_58_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_58_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_58_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_58_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_58_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_58_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_58_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_58_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_59_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_59_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_59_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_59_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_59_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_59_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_59_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_59_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_59_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_59_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_60_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_60_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_60_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_60_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_60_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_60_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_60_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_60_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_60_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_60_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_61_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_61_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_61_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_61_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_61_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_61_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_61_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_61_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_61_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_61_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_62_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_62_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_62_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_62_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_62_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_62_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_62_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_62_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_62_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_62_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_63_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_63_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_63_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_63_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_63_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_63_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_63_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_63_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_63_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_63_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_64_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_64_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_64_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_64_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_64_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_64_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_64_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_64_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_64_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_64_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_65_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_65_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_65_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_65_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_65_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_65_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_65_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_65_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_65_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_65_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_66_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_66_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_66_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_66_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_66_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_66_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_66_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_66_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_66_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_66_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_67_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_67_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_67_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_67_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_67_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_67_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_67_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_67_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_67_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_67_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_68_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_68_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_68_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_68_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_68_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_68_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_68_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_68_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_68_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_68_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_69_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_69_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_69_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_69_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_69_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_69_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_69_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_69_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_69_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_69_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_70_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_70_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_70_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_70_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_70_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_70_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_70_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_70_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_70_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_70_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_71_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_71_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_71_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_71_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_71_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_71_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_71_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_71_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_71_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_71_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_72_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_72_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_72_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_72_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_72_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_72_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_72_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_72_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_72_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_72_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_73_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_73_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_73_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_73_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_73_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_73_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_73_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_73_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_73_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_73_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_74_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_74_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_74_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_74_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_74_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_74_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_74_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_74_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_74_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_74_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_75_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_75_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_75_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_75_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_75_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_75_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_75_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_75_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_75_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_75_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_76_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_76_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_76_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_76_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_76_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_76_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_76_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_76_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_76_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_76_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_77_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_77_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_77_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_77_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_77_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_77_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_77_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_77_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_77_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_77_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_78_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_78_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_78_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_78_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_78_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_78_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_78_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_78_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_78_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_78_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_79_clock; // @[FFTDesigns.scala 3122:34]
  wire  DFT_r_v2_79_reset; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_79_io_in_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_79_io_in_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_79_io_in_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_79_io_in_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_79_io_out_0_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_79_io_out_0_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_79_io_out_1_Re; // @[FFTDesigns.scala 3122:34]
  wire [31:0] DFT_r_v2_79_io_out_1_Im; // @[FFTDesigns.scala 3122:34]
  wire [31:0] PermutationsBasic_io_in_0_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_0_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_1_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_1_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_2_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_2_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_3_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_3_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_4_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_4_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_5_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_5_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_6_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_6_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_7_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_7_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_8_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_8_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_9_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_9_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_10_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_10_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_11_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_11_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_12_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_12_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_13_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_13_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_14_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_14_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_15_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_15_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_16_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_16_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_17_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_17_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_18_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_18_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_19_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_19_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_20_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_20_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_21_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_21_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_22_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_22_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_23_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_23_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_24_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_24_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_25_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_25_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_26_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_26_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_27_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_27_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_28_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_28_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_29_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_29_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_30_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_30_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_31_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_in_31_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_0_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_0_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_1_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_1_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_2_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_2_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_3_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_3_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_4_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_4_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_5_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_5_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_6_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_6_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_7_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_7_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_8_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_8_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_9_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_9_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_10_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_10_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_11_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_11_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_12_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_12_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_13_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_13_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_14_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_14_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_15_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_15_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_16_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_16_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_17_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_17_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_18_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_18_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_19_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_19_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_20_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_20_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_21_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_21_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_22_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_22_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_23_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_23_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_24_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_24_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_25_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_25_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_26_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_26_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_27_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_27_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_28_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_28_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_29_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_29_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_30_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_30_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_31_Re; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_io_out_31_Im; // @[FFTDesigns.scala 3127:35]
  wire [31:0] PermutationsBasic_1_io_in_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_in_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_1_io_out_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_in_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_2_io_out_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_in_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_3_io_out_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_in_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_4_io_out_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_in_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_0_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_0_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_1_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_1_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_2_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_2_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_3_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_3_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_4_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_4_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_5_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_5_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_6_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_6_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_7_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_7_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_8_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_8_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_9_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_9_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_10_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_10_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_11_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_11_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_12_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_12_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_13_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_13_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_14_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_14_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_15_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_15_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_16_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_16_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_17_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_17_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_18_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_18_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_19_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_19_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_20_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_20_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_21_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_21_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_22_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_22_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_23_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_23_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_24_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_24_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_25_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_25_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_26_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_26_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_27_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_27_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_28_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_28_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_29_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_29_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_30_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_30_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_31_Re; // @[FFTDesigns.scala 3129:37]
  wire [31:0] PermutationsBasic_5_io_out_31_Im; // @[FFTDesigns.scala 3129:37]
  wire [31:0] TwiddleFactors_io_in_0_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_0_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_1_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_1_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_2_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_2_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_3_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_3_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_4_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_4_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_5_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_5_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_6_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_6_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_7_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_7_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_8_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_8_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_9_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_9_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_10_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_10_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_11_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_11_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_12_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_12_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_13_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_13_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_14_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_14_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_15_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_15_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_16_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_16_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_17_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_17_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_18_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_18_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_19_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_19_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_20_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_20_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_21_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_21_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_22_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_22_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_23_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_23_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_24_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_24_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_25_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_25_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_26_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_26_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_27_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_27_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_28_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_28_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_29_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_29_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_30_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_30_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_31_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_in_31_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_0_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_0_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_1_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_1_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_2_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_2_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_3_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_3_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_4_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_4_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_5_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_5_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_6_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_6_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_7_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_7_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_8_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_8_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_9_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_9_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_10_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_10_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_11_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_11_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_12_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_12_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_13_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_13_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_14_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_14_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_15_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_15_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_16_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_16_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_17_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_17_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_18_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_18_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_19_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_19_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_20_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_20_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_21_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_21_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_22_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_22_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_23_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_23_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_24_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_24_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_25_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_25_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_26_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_26_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_27_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_27_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_28_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_28_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_29_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_29_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_30_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_30_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_31_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_io_out_31_Im; // @[FFTDesigns.scala 3133:24]
  wire  TwiddleFactors_1_clock; // @[FFTDesigns.scala 3133:24]
  wire  TwiddleFactors_1_reset; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_0_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_0_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_1_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_1_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_2_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_2_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_3_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_3_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_4_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_4_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_5_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_5_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_6_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_6_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_7_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_7_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_8_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_8_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_9_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_9_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_10_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_10_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_11_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_11_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_12_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_12_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_13_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_13_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_14_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_14_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_15_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_15_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_16_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_16_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_17_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_17_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_18_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_18_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_19_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_19_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_20_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_20_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_21_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_21_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_22_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_22_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_23_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_23_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_24_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_24_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_25_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_25_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_26_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_26_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_27_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_27_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_28_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_28_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_29_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_29_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_30_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_30_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_31_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_in_31_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_0_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_0_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_1_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_1_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_2_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_2_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_3_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_3_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_4_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_4_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_5_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_5_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_6_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_6_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_7_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_7_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_8_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_8_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_9_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_9_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_10_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_10_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_11_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_11_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_12_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_12_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_13_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_13_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_14_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_14_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_15_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_15_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_16_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_16_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_17_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_17_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_18_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_18_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_19_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_19_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_20_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_20_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_21_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_21_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_22_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_22_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_23_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_23_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_24_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_24_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_25_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_25_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_26_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_26_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_27_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_27_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_28_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_28_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_29_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_29_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_30_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_30_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_31_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_1_io_out_31_Im; // @[FFTDesigns.scala 3133:24]
  wire  TwiddleFactors_2_clock; // @[FFTDesigns.scala 3133:24]
  wire  TwiddleFactors_2_reset; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_0_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_0_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_1_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_1_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_2_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_2_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_3_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_3_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_4_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_4_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_5_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_5_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_6_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_6_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_7_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_7_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_8_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_8_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_9_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_9_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_10_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_10_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_11_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_11_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_12_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_12_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_13_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_13_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_14_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_14_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_15_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_15_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_16_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_16_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_17_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_17_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_18_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_18_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_19_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_19_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_20_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_20_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_21_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_21_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_22_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_22_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_23_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_23_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_24_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_24_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_25_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_25_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_26_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_26_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_27_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_27_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_28_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_28_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_29_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_29_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_30_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_30_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_31_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_in_31_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_0_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_0_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_1_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_1_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_2_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_2_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_3_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_3_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_4_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_4_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_5_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_5_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_6_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_6_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_7_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_7_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_8_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_8_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_9_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_9_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_10_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_10_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_11_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_11_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_12_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_12_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_13_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_13_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_14_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_14_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_15_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_15_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_16_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_16_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_17_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_17_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_18_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_18_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_19_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_19_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_20_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_20_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_21_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_21_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_22_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_22_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_23_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_23_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_24_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_24_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_25_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_25_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_26_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_26_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_27_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_27_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_28_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_28_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_29_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_29_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_30_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_30_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_31_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_2_io_out_31_Im; // @[FFTDesigns.scala 3133:24]
  wire  TwiddleFactors_3_clock; // @[FFTDesigns.scala 3133:24]
  wire  TwiddleFactors_3_reset; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_0_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_0_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_1_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_1_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_2_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_2_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_3_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_3_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_4_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_4_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_5_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_5_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_6_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_6_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_7_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_7_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_8_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_8_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_9_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_9_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_10_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_10_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_11_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_11_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_12_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_12_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_13_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_13_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_14_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_14_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_15_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_15_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_16_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_16_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_17_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_17_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_18_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_18_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_19_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_19_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_20_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_20_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_21_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_21_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_22_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_22_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_23_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_23_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_24_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_24_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_25_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_25_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_26_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_26_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_27_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_27_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_28_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_28_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_29_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_29_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_30_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_30_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_31_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_in_31_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_0_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_0_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_1_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_1_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_2_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_2_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_3_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_3_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_4_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_4_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_5_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_5_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_6_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_6_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_7_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_7_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_8_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_8_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_9_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_9_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_10_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_10_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_11_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_11_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_12_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_12_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_13_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_13_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_14_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_14_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_15_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_15_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_16_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_16_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_17_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_17_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_18_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_18_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_19_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_19_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_20_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_20_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_21_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_21_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_22_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_22_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_23_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_23_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_24_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_24_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_25_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_25_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_26_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_26_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_27_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_27_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_28_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_28_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_29_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_29_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_30_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_30_Im; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_31_Re; // @[FFTDesigns.scala 3133:24]
  wire [31:0] TwiddleFactors_3_io_out_31_Im; // @[FFTDesigns.scala 3133:24]
  DFT_r_v2_32 DFT_r_v2 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_clock),
    .reset(DFT_r_v2_reset),
    .io_in_0_Re(DFT_r_v2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_1 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_1_clock),
    .reset(DFT_r_v2_1_reset),
    .io_in_0_Re(DFT_r_v2_1_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_1_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_1_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_1_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_1_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_1_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_1_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_1_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_2 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_2_clock),
    .reset(DFT_r_v2_2_reset),
    .io_in_0_Re(DFT_r_v2_2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_2_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_2_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_3 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_3_clock),
    .reset(DFT_r_v2_3_reset),
    .io_in_0_Re(DFT_r_v2_3_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_3_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_3_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_3_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_3_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_3_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_3_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_3_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_4 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_4_clock),
    .reset(DFT_r_v2_4_reset),
    .io_in_0_Re(DFT_r_v2_4_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_4_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_4_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_4_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_4_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_4_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_4_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_4_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_5 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_5_clock),
    .reset(DFT_r_v2_5_reset),
    .io_in_0_Re(DFT_r_v2_5_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_5_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_5_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_5_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_5_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_5_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_5_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_5_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_6 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_6_clock),
    .reset(DFT_r_v2_6_reset),
    .io_in_0_Re(DFT_r_v2_6_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_6_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_6_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_6_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_6_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_6_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_6_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_6_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_7 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_7_clock),
    .reset(DFT_r_v2_7_reset),
    .io_in_0_Re(DFT_r_v2_7_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_7_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_7_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_7_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_7_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_7_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_7_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_7_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_8 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_8_clock),
    .reset(DFT_r_v2_8_reset),
    .io_in_0_Re(DFT_r_v2_8_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_8_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_8_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_8_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_8_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_8_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_8_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_8_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_9 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_9_clock),
    .reset(DFT_r_v2_9_reset),
    .io_in_0_Re(DFT_r_v2_9_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_9_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_9_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_9_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_9_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_9_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_9_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_9_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_10 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_10_clock),
    .reset(DFT_r_v2_10_reset),
    .io_in_0_Re(DFT_r_v2_10_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_10_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_10_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_10_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_10_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_10_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_10_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_10_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_11 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_11_clock),
    .reset(DFT_r_v2_11_reset),
    .io_in_0_Re(DFT_r_v2_11_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_11_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_11_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_11_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_11_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_11_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_11_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_11_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_12 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_12_clock),
    .reset(DFT_r_v2_12_reset),
    .io_in_0_Re(DFT_r_v2_12_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_12_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_12_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_12_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_12_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_12_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_12_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_12_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_13 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_13_clock),
    .reset(DFT_r_v2_13_reset),
    .io_in_0_Re(DFT_r_v2_13_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_13_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_13_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_13_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_13_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_13_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_13_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_13_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_14 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_14_clock),
    .reset(DFT_r_v2_14_reset),
    .io_in_0_Re(DFT_r_v2_14_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_14_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_14_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_14_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_14_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_14_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_14_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_14_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_15 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_15_clock),
    .reset(DFT_r_v2_15_reset),
    .io_in_0_Re(DFT_r_v2_15_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_15_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_15_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_15_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_15_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_15_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_15_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_15_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_16 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_16_clock),
    .reset(DFT_r_v2_16_reset),
    .io_in_0_Re(DFT_r_v2_16_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_16_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_16_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_16_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_16_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_16_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_16_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_16_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_17 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_17_clock),
    .reset(DFT_r_v2_17_reset),
    .io_in_0_Re(DFT_r_v2_17_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_17_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_17_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_17_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_17_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_17_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_17_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_17_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_18 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_18_clock),
    .reset(DFT_r_v2_18_reset),
    .io_in_0_Re(DFT_r_v2_18_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_18_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_18_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_18_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_18_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_18_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_18_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_18_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_19 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_19_clock),
    .reset(DFT_r_v2_19_reset),
    .io_in_0_Re(DFT_r_v2_19_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_19_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_19_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_19_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_19_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_19_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_19_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_19_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_20 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_20_clock),
    .reset(DFT_r_v2_20_reset),
    .io_in_0_Re(DFT_r_v2_20_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_20_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_20_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_20_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_20_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_20_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_20_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_20_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_21 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_21_clock),
    .reset(DFT_r_v2_21_reset),
    .io_in_0_Re(DFT_r_v2_21_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_21_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_21_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_21_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_21_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_21_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_21_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_21_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_22 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_22_clock),
    .reset(DFT_r_v2_22_reset),
    .io_in_0_Re(DFT_r_v2_22_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_22_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_22_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_22_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_22_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_22_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_22_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_22_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_23 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_23_clock),
    .reset(DFT_r_v2_23_reset),
    .io_in_0_Re(DFT_r_v2_23_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_23_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_23_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_23_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_23_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_23_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_23_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_23_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_24 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_24_clock),
    .reset(DFT_r_v2_24_reset),
    .io_in_0_Re(DFT_r_v2_24_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_24_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_24_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_24_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_24_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_24_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_24_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_24_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_25 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_25_clock),
    .reset(DFT_r_v2_25_reset),
    .io_in_0_Re(DFT_r_v2_25_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_25_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_25_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_25_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_25_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_25_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_25_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_25_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_26 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_26_clock),
    .reset(DFT_r_v2_26_reset),
    .io_in_0_Re(DFT_r_v2_26_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_26_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_26_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_26_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_26_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_26_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_26_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_26_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_27 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_27_clock),
    .reset(DFT_r_v2_27_reset),
    .io_in_0_Re(DFT_r_v2_27_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_27_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_27_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_27_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_27_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_27_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_27_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_27_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_28 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_28_clock),
    .reset(DFT_r_v2_28_reset),
    .io_in_0_Re(DFT_r_v2_28_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_28_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_28_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_28_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_28_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_28_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_28_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_28_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_29 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_29_clock),
    .reset(DFT_r_v2_29_reset),
    .io_in_0_Re(DFT_r_v2_29_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_29_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_29_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_29_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_29_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_29_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_29_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_29_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_30 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_30_clock),
    .reset(DFT_r_v2_30_reset),
    .io_in_0_Re(DFT_r_v2_30_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_30_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_30_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_30_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_30_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_30_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_30_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_30_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_31 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_31_clock),
    .reset(DFT_r_v2_31_reset),
    .io_in_0_Re(DFT_r_v2_31_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_31_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_31_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_31_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_31_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_31_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_31_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_31_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_32 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_32_clock),
    .reset(DFT_r_v2_32_reset),
    .io_in_0_Re(DFT_r_v2_32_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_32_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_32_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_32_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_32_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_32_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_32_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_32_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_33 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_33_clock),
    .reset(DFT_r_v2_33_reset),
    .io_in_0_Re(DFT_r_v2_33_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_33_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_33_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_33_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_33_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_33_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_33_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_33_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_34 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_34_clock),
    .reset(DFT_r_v2_34_reset),
    .io_in_0_Re(DFT_r_v2_34_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_34_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_34_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_34_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_34_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_34_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_34_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_34_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_35 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_35_clock),
    .reset(DFT_r_v2_35_reset),
    .io_in_0_Re(DFT_r_v2_35_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_35_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_35_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_35_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_35_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_35_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_35_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_35_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_36 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_36_clock),
    .reset(DFT_r_v2_36_reset),
    .io_in_0_Re(DFT_r_v2_36_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_36_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_36_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_36_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_36_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_36_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_36_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_36_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_37 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_37_clock),
    .reset(DFT_r_v2_37_reset),
    .io_in_0_Re(DFT_r_v2_37_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_37_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_37_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_37_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_37_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_37_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_37_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_37_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_38 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_38_clock),
    .reset(DFT_r_v2_38_reset),
    .io_in_0_Re(DFT_r_v2_38_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_38_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_38_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_38_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_38_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_38_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_38_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_38_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_39 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_39_clock),
    .reset(DFT_r_v2_39_reset),
    .io_in_0_Re(DFT_r_v2_39_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_39_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_39_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_39_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_39_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_39_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_39_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_39_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_40 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_40_clock),
    .reset(DFT_r_v2_40_reset),
    .io_in_0_Re(DFT_r_v2_40_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_40_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_40_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_40_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_40_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_40_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_40_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_40_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_41 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_41_clock),
    .reset(DFT_r_v2_41_reset),
    .io_in_0_Re(DFT_r_v2_41_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_41_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_41_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_41_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_41_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_41_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_41_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_41_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_42 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_42_clock),
    .reset(DFT_r_v2_42_reset),
    .io_in_0_Re(DFT_r_v2_42_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_42_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_42_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_42_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_42_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_42_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_42_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_42_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_43 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_43_clock),
    .reset(DFT_r_v2_43_reset),
    .io_in_0_Re(DFT_r_v2_43_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_43_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_43_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_43_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_43_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_43_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_43_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_43_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_44 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_44_clock),
    .reset(DFT_r_v2_44_reset),
    .io_in_0_Re(DFT_r_v2_44_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_44_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_44_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_44_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_44_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_44_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_44_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_44_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_45 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_45_clock),
    .reset(DFT_r_v2_45_reset),
    .io_in_0_Re(DFT_r_v2_45_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_45_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_45_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_45_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_45_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_45_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_45_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_45_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_46 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_46_clock),
    .reset(DFT_r_v2_46_reset),
    .io_in_0_Re(DFT_r_v2_46_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_46_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_46_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_46_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_46_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_46_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_46_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_46_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_47 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_47_clock),
    .reset(DFT_r_v2_47_reset),
    .io_in_0_Re(DFT_r_v2_47_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_47_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_47_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_47_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_47_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_47_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_47_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_47_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_48 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_48_clock),
    .reset(DFT_r_v2_48_reset),
    .io_in_0_Re(DFT_r_v2_48_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_48_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_48_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_48_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_48_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_48_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_48_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_48_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_49 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_49_clock),
    .reset(DFT_r_v2_49_reset),
    .io_in_0_Re(DFT_r_v2_49_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_49_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_49_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_49_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_49_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_49_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_49_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_49_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_50 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_50_clock),
    .reset(DFT_r_v2_50_reset),
    .io_in_0_Re(DFT_r_v2_50_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_50_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_50_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_50_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_50_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_50_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_50_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_50_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_51 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_51_clock),
    .reset(DFT_r_v2_51_reset),
    .io_in_0_Re(DFT_r_v2_51_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_51_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_51_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_51_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_51_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_51_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_51_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_51_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_52 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_52_clock),
    .reset(DFT_r_v2_52_reset),
    .io_in_0_Re(DFT_r_v2_52_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_52_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_52_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_52_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_52_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_52_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_52_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_52_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_53 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_53_clock),
    .reset(DFT_r_v2_53_reset),
    .io_in_0_Re(DFT_r_v2_53_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_53_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_53_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_53_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_53_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_53_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_53_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_53_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_54 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_54_clock),
    .reset(DFT_r_v2_54_reset),
    .io_in_0_Re(DFT_r_v2_54_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_54_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_54_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_54_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_54_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_54_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_54_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_54_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_55 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_55_clock),
    .reset(DFT_r_v2_55_reset),
    .io_in_0_Re(DFT_r_v2_55_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_55_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_55_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_55_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_55_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_55_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_55_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_55_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_56 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_56_clock),
    .reset(DFT_r_v2_56_reset),
    .io_in_0_Re(DFT_r_v2_56_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_56_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_56_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_56_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_56_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_56_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_56_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_56_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_57 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_57_clock),
    .reset(DFT_r_v2_57_reset),
    .io_in_0_Re(DFT_r_v2_57_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_57_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_57_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_57_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_57_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_57_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_57_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_57_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_58 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_58_clock),
    .reset(DFT_r_v2_58_reset),
    .io_in_0_Re(DFT_r_v2_58_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_58_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_58_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_58_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_58_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_58_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_58_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_58_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_59 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_59_clock),
    .reset(DFT_r_v2_59_reset),
    .io_in_0_Re(DFT_r_v2_59_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_59_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_59_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_59_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_59_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_59_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_59_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_59_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_60 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_60_clock),
    .reset(DFT_r_v2_60_reset),
    .io_in_0_Re(DFT_r_v2_60_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_60_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_60_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_60_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_60_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_60_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_60_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_60_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_61 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_61_clock),
    .reset(DFT_r_v2_61_reset),
    .io_in_0_Re(DFT_r_v2_61_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_61_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_61_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_61_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_61_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_61_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_61_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_61_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_62 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_62_clock),
    .reset(DFT_r_v2_62_reset),
    .io_in_0_Re(DFT_r_v2_62_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_62_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_62_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_62_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_62_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_62_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_62_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_62_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_63 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_63_clock),
    .reset(DFT_r_v2_63_reset),
    .io_in_0_Re(DFT_r_v2_63_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_63_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_63_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_63_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_63_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_63_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_63_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_63_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_64 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_64_clock),
    .reset(DFT_r_v2_64_reset),
    .io_in_0_Re(DFT_r_v2_64_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_64_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_64_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_64_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_64_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_64_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_64_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_64_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_65 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_65_clock),
    .reset(DFT_r_v2_65_reset),
    .io_in_0_Re(DFT_r_v2_65_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_65_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_65_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_65_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_65_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_65_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_65_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_65_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_66 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_66_clock),
    .reset(DFT_r_v2_66_reset),
    .io_in_0_Re(DFT_r_v2_66_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_66_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_66_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_66_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_66_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_66_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_66_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_66_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_67 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_67_clock),
    .reset(DFT_r_v2_67_reset),
    .io_in_0_Re(DFT_r_v2_67_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_67_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_67_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_67_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_67_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_67_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_67_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_67_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_68 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_68_clock),
    .reset(DFT_r_v2_68_reset),
    .io_in_0_Re(DFT_r_v2_68_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_68_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_68_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_68_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_68_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_68_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_68_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_68_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_69 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_69_clock),
    .reset(DFT_r_v2_69_reset),
    .io_in_0_Re(DFT_r_v2_69_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_69_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_69_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_69_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_69_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_69_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_69_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_69_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_70 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_70_clock),
    .reset(DFT_r_v2_70_reset),
    .io_in_0_Re(DFT_r_v2_70_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_70_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_70_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_70_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_70_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_70_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_70_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_70_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_71 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_71_clock),
    .reset(DFT_r_v2_71_reset),
    .io_in_0_Re(DFT_r_v2_71_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_71_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_71_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_71_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_71_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_71_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_71_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_71_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_72 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_72_clock),
    .reset(DFT_r_v2_72_reset),
    .io_in_0_Re(DFT_r_v2_72_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_72_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_72_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_72_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_72_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_72_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_72_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_72_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_73 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_73_clock),
    .reset(DFT_r_v2_73_reset),
    .io_in_0_Re(DFT_r_v2_73_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_73_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_73_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_73_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_73_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_73_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_73_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_73_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_74 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_74_clock),
    .reset(DFT_r_v2_74_reset),
    .io_in_0_Re(DFT_r_v2_74_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_74_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_74_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_74_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_74_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_74_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_74_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_74_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_75 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_75_clock),
    .reset(DFT_r_v2_75_reset),
    .io_in_0_Re(DFT_r_v2_75_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_75_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_75_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_75_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_75_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_75_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_75_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_75_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_76 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_76_clock),
    .reset(DFT_r_v2_76_reset),
    .io_in_0_Re(DFT_r_v2_76_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_76_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_76_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_76_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_76_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_76_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_76_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_76_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_77 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_77_clock),
    .reset(DFT_r_v2_77_reset),
    .io_in_0_Re(DFT_r_v2_77_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_77_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_77_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_77_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_77_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_77_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_77_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_77_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_78 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_78_clock),
    .reset(DFT_r_v2_78_reset),
    .io_in_0_Re(DFT_r_v2_78_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_78_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_78_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_78_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_78_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_78_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_78_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_78_io_out_1_Im)
  );
  DFT_r_v2_32 DFT_r_v2_79 ( // @[FFTDesigns.scala 3122:34]
    .clock(DFT_r_v2_79_clock),
    .reset(DFT_r_v2_79_reset),
    .io_in_0_Re(DFT_r_v2_79_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_79_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_79_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_79_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_79_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_79_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_79_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_79_io_out_1_Im)
  );
  PermutationsBasic_64 PermutationsBasic ( // @[FFTDesigns.scala 3127:35]
    .io_in_0_Re(PermutationsBasic_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_io_in_31_Im),
    .io_out_0_Re(PermutationsBasic_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_io_out_31_Im)
  );
  PermutationsBasic_65 PermutationsBasic_1 ( // @[FFTDesigns.scala 3129:37]
    .io_in_0_Re(PermutationsBasic_1_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_1_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_1_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_1_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_1_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_1_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_1_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_1_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_1_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_1_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_1_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_1_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_1_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_1_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_1_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_1_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_1_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_1_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_1_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_1_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_1_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_1_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_1_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_1_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_1_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_1_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_1_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_1_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_1_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_1_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_1_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_1_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_1_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_1_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_1_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_1_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_1_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_1_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_1_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_1_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_1_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_1_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_1_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_1_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_1_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_1_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_1_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_1_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_1_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_1_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_1_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_1_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_1_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_1_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_1_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_1_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_1_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_1_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_1_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_1_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_1_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_1_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_1_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_1_io_in_31_Im),
    .io_out_0_Re(PermutationsBasic_1_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_1_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_1_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_1_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_1_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_1_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_1_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_1_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_1_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_1_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_1_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_1_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_1_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_1_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_1_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_1_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_1_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_1_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_1_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_1_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_1_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_1_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_1_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_1_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_1_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_1_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_1_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_1_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_1_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_1_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_1_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_1_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_1_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_1_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_1_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_1_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_1_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_1_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_1_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_1_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_1_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_1_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_1_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_1_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_1_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_1_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_1_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_1_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_1_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_1_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_1_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_1_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_1_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_1_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_1_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_1_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_1_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_1_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_1_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_1_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_1_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_1_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_1_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_1_io_out_31_Im)
  );
  PermutationsBasic_65 PermutationsBasic_2 ( // @[FFTDesigns.scala 3129:37]
    .io_in_0_Re(PermutationsBasic_2_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_2_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_2_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_2_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_2_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_2_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_2_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_2_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_2_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_2_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_2_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_2_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_2_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_2_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_2_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_2_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_2_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_2_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_2_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_2_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_2_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_2_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_2_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_2_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_2_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_2_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_2_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_2_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_2_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_2_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_2_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_2_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_2_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_2_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_2_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_2_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_2_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_2_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_2_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_2_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_2_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_2_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_2_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_2_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_2_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_2_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_2_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_2_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_2_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_2_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_2_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_2_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_2_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_2_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_2_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_2_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_2_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_2_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_2_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_2_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_2_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_2_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_2_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_2_io_in_31_Im),
    .io_out_0_Re(PermutationsBasic_2_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_2_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_2_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_2_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_2_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_2_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_2_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_2_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_2_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_2_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_2_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_2_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_2_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_2_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_2_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_2_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_2_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_2_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_2_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_2_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_2_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_2_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_2_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_2_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_2_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_2_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_2_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_2_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_2_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_2_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_2_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_2_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_2_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_2_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_2_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_2_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_2_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_2_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_2_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_2_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_2_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_2_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_2_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_2_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_2_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_2_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_2_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_2_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_2_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_2_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_2_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_2_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_2_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_2_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_2_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_2_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_2_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_2_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_2_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_2_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_2_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_2_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_2_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_2_io_out_31_Im)
  );
  PermutationsBasic_65 PermutationsBasic_3 ( // @[FFTDesigns.scala 3129:37]
    .io_in_0_Re(PermutationsBasic_3_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_3_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_3_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_3_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_3_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_3_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_3_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_3_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_3_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_3_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_3_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_3_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_3_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_3_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_3_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_3_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_3_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_3_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_3_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_3_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_3_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_3_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_3_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_3_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_3_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_3_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_3_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_3_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_3_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_3_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_3_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_3_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_3_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_3_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_3_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_3_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_3_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_3_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_3_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_3_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_3_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_3_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_3_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_3_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_3_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_3_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_3_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_3_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_3_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_3_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_3_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_3_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_3_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_3_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_3_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_3_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_3_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_3_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_3_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_3_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_3_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_3_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_3_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_3_io_in_31_Im),
    .io_out_0_Re(PermutationsBasic_3_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_3_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_3_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_3_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_3_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_3_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_3_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_3_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_3_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_3_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_3_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_3_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_3_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_3_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_3_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_3_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_3_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_3_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_3_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_3_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_3_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_3_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_3_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_3_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_3_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_3_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_3_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_3_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_3_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_3_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_3_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_3_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_3_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_3_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_3_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_3_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_3_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_3_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_3_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_3_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_3_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_3_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_3_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_3_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_3_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_3_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_3_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_3_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_3_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_3_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_3_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_3_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_3_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_3_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_3_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_3_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_3_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_3_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_3_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_3_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_3_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_3_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_3_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_3_io_out_31_Im)
  );
  PermutationsBasic_65 PermutationsBasic_4 ( // @[FFTDesigns.scala 3129:37]
    .io_in_0_Re(PermutationsBasic_4_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_4_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_4_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_4_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_4_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_4_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_4_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_4_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_4_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_4_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_4_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_4_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_4_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_4_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_4_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_4_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_4_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_4_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_4_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_4_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_4_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_4_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_4_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_4_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_4_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_4_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_4_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_4_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_4_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_4_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_4_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_4_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_4_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_4_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_4_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_4_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_4_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_4_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_4_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_4_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_4_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_4_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_4_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_4_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_4_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_4_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_4_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_4_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_4_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_4_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_4_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_4_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_4_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_4_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_4_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_4_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_4_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_4_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_4_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_4_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_4_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_4_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_4_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_4_io_in_31_Im),
    .io_out_0_Re(PermutationsBasic_4_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_4_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_4_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_4_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_4_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_4_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_4_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_4_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_4_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_4_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_4_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_4_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_4_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_4_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_4_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_4_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_4_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_4_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_4_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_4_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_4_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_4_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_4_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_4_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_4_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_4_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_4_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_4_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_4_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_4_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_4_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_4_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_4_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_4_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_4_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_4_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_4_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_4_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_4_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_4_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_4_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_4_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_4_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_4_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_4_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_4_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_4_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_4_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_4_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_4_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_4_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_4_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_4_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_4_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_4_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_4_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_4_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_4_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_4_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_4_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_4_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_4_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_4_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_4_io_out_31_Im)
  );
  PermutationsBasic_65 PermutationsBasic_5 ( // @[FFTDesigns.scala 3129:37]
    .io_in_0_Re(PermutationsBasic_5_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_5_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_5_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_5_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_5_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_5_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_5_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_5_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_5_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_5_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_5_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_5_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_5_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_5_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_5_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_5_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_5_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_5_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_5_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_5_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_5_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_5_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_5_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_5_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_5_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_5_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_5_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_5_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_5_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_5_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_5_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_5_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_5_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_5_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_5_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_5_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_5_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_5_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_5_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_5_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_5_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_5_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_5_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_5_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_5_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_5_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_5_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_5_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_5_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_5_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_5_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_5_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_5_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_5_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_5_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_5_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_5_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_5_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_5_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_5_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_5_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_5_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_5_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_5_io_in_31_Im),
    .io_out_0_Re(PermutationsBasic_5_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_5_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_5_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_5_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_5_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_5_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_5_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_5_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_5_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_5_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_5_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_5_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_5_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_5_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_5_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_5_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_5_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_5_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_5_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_5_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_5_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_5_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_5_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_5_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_5_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_5_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_5_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_5_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_5_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_5_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_5_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_5_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_5_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_5_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_5_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_5_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_5_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_5_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_5_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_5_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_5_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_5_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_5_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_5_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_5_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_5_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_5_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_5_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_5_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_5_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_5_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_5_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_5_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_5_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_5_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_5_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_5_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_5_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_5_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_5_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_5_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_5_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_5_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_5_io_out_31_Im)
  );
  TwiddleFactors TwiddleFactors ( // @[FFTDesigns.scala 3133:24]
    .io_in_0_Re(TwiddleFactors_io_in_0_Re),
    .io_in_0_Im(TwiddleFactors_io_in_0_Im),
    .io_in_1_Re(TwiddleFactors_io_in_1_Re),
    .io_in_1_Im(TwiddleFactors_io_in_1_Im),
    .io_in_2_Re(TwiddleFactors_io_in_2_Re),
    .io_in_2_Im(TwiddleFactors_io_in_2_Im),
    .io_in_3_Re(TwiddleFactors_io_in_3_Re),
    .io_in_3_Im(TwiddleFactors_io_in_3_Im),
    .io_in_4_Re(TwiddleFactors_io_in_4_Re),
    .io_in_4_Im(TwiddleFactors_io_in_4_Im),
    .io_in_5_Re(TwiddleFactors_io_in_5_Re),
    .io_in_5_Im(TwiddleFactors_io_in_5_Im),
    .io_in_6_Re(TwiddleFactors_io_in_6_Re),
    .io_in_6_Im(TwiddleFactors_io_in_6_Im),
    .io_in_7_Re(TwiddleFactors_io_in_7_Re),
    .io_in_7_Im(TwiddleFactors_io_in_7_Im),
    .io_in_8_Re(TwiddleFactors_io_in_8_Re),
    .io_in_8_Im(TwiddleFactors_io_in_8_Im),
    .io_in_9_Re(TwiddleFactors_io_in_9_Re),
    .io_in_9_Im(TwiddleFactors_io_in_9_Im),
    .io_in_10_Re(TwiddleFactors_io_in_10_Re),
    .io_in_10_Im(TwiddleFactors_io_in_10_Im),
    .io_in_11_Re(TwiddleFactors_io_in_11_Re),
    .io_in_11_Im(TwiddleFactors_io_in_11_Im),
    .io_in_12_Re(TwiddleFactors_io_in_12_Re),
    .io_in_12_Im(TwiddleFactors_io_in_12_Im),
    .io_in_13_Re(TwiddleFactors_io_in_13_Re),
    .io_in_13_Im(TwiddleFactors_io_in_13_Im),
    .io_in_14_Re(TwiddleFactors_io_in_14_Re),
    .io_in_14_Im(TwiddleFactors_io_in_14_Im),
    .io_in_15_Re(TwiddleFactors_io_in_15_Re),
    .io_in_15_Im(TwiddleFactors_io_in_15_Im),
    .io_in_16_Re(TwiddleFactors_io_in_16_Re),
    .io_in_16_Im(TwiddleFactors_io_in_16_Im),
    .io_in_17_Re(TwiddleFactors_io_in_17_Re),
    .io_in_17_Im(TwiddleFactors_io_in_17_Im),
    .io_in_18_Re(TwiddleFactors_io_in_18_Re),
    .io_in_18_Im(TwiddleFactors_io_in_18_Im),
    .io_in_19_Re(TwiddleFactors_io_in_19_Re),
    .io_in_19_Im(TwiddleFactors_io_in_19_Im),
    .io_in_20_Re(TwiddleFactors_io_in_20_Re),
    .io_in_20_Im(TwiddleFactors_io_in_20_Im),
    .io_in_21_Re(TwiddleFactors_io_in_21_Re),
    .io_in_21_Im(TwiddleFactors_io_in_21_Im),
    .io_in_22_Re(TwiddleFactors_io_in_22_Re),
    .io_in_22_Im(TwiddleFactors_io_in_22_Im),
    .io_in_23_Re(TwiddleFactors_io_in_23_Re),
    .io_in_23_Im(TwiddleFactors_io_in_23_Im),
    .io_in_24_Re(TwiddleFactors_io_in_24_Re),
    .io_in_24_Im(TwiddleFactors_io_in_24_Im),
    .io_in_25_Re(TwiddleFactors_io_in_25_Re),
    .io_in_25_Im(TwiddleFactors_io_in_25_Im),
    .io_in_26_Re(TwiddleFactors_io_in_26_Re),
    .io_in_26_Im(TwiddleFactors_io_in_26_Im),
    .io_in_27_Re(TwiddleFactors_io_in_27_Re),
    .io_in_27_Im(TwiddleFactors_io_in_27_Im),
    .io_in_28_Re(TwiddleFactors_io_in_28_Re),
    .io_in_28_Im(TwiddleFactors_io_in_28_Im),
    .io_in_29_Re(TwiddleFactors_io_in_29_Re),
    .io_in_29_Im(TwiddleFactors_io_in_29_Im),
    .io_in_30_Re(TwiddleFactors_io_in_30_Re),
    .io_in_30_Im(TwiddleFactors_io_in_30_Im),
    .io_in_31_Re(TwiddleFactors_io_in_31_Re),
    .io_in_31_Im(TwiddleFactors_io_in_31_Im),
    .io_out_0_Re(TwiddleFactors_io_out_0_Re),
    .io_out_0_Im(TwiddleFactors_io_out_0_Im),
    .io_out_1_Re(TwiddleFactors_io_out_1_Re),
    .io_out_1_Im(TwiddleFactors_io_out_1_Im),
    .io_out_2_Re(TwiddleFactors_io_out_2_Re),
    .io_out_2_Im(TwiddleFactors_io_out_2_Im),
    .io_out_3_Re(TwiddleFactors_io_out_3_Re),
    .io_out_3_Im(TwiddleFactors_io_out_3_Im),
    .io_out_4_Re(TwiddleFactors_io_out_4_Re),
    .io_out_4_Im(TwiddleFactors_io_out_4_Im),
    .io_out_5_Re(TwiddleFactors_io_out_5_Re),
    .io_out_5_Im(TwiddleFactors_io_out_5_Im),
    .io_out_6_Re(TwiddleFactors_io_out_6_Re),
    .io_out_6_Im(TwiddleFactors_io_out_6_Im),
    .io_out_7_Re(TwiddleFactors_io_out_7_Re),
    .io_out_7_Im(TwiddleFactors_io_out_7_Im),
    .io_out_8_Re(TwiddleFactors_io_out_8_Re),
    .io_out_8_Im(TwiddleFactors_io_out_8_Im),
    .io_out_9_Re(TwiddleFactors_io_out_9_Re),
    .io_out_9_Im(TwiddleFactors_io_out_9_Im),
    .io_out_10_Re(TwiddleFactors_io_out_10_Re),
    .io_out_10_Im(TwiddleFactors_io_out_10_Im),
    .io_out_11_Re(TwiddleFactors_io_out_11_Re),
    .io_out_11_Im(TwiddleFactors_io_out_11_Im),
    .io_out_12_Re(TwiddleFactors_io_out_12_Re),
    .io_out_12_Im(TwiddleFactors_io_out_12_Im),
    .io_out_13_Re(TwiddleFactors_io_out_13_Re),
    .io_out_13_Im(TwiddleFactors_io_out_13_Im),
    .io_out_14_Re(TwiddleFactors_io_out_14_Re),
    .io_out_14_Im(TwiddleFactors_io_out_14_Im),
    .io_out_15_Re(TwiddleFactors_io_out_15_Re),
    .io_out_15_Im(TwiddleFactors_io_out_15_Im),
    .io_out_16_Re(TwiddleFactors_io_out_16_Re),
    .io_out_16_Im(TwiddleFactors_io_out_16_Im),
    .io_out_17_Re(TwiddleFactors_io_out_17_Re),
    .io_out_17_Im(TwiddleFactors_io_out_17_Im),
    .io_out_18_Re(TwiddleFactors_io_out_18_Re),
    .io_out_18_Im(TwiddleFactors_io_out_18_Im),
    .io_out_19_Re(TwiddleFactors_io_out_19_Re),
    .io_out_19_Im(TwiddleFactors_io_out_19_Im),
    .io_out_20_Re(TwiddleFactors_io_out_20_Re),
    .io_out_20_Im(TwiddleFactors_io_out_20_Im),
    .io_out_21_Re(TwiddleFactors_io_out_21_Re),
    .io_out_21_Im(TwiddleFactors_io_out_21_Im),
    .io_out_22_Re(TwiddleFactors_io_out_22_Re),
    .io_out_22_Im(TwiddleFactors_io_out_22_Im),
    .io_out_23_Re(TwiddleFactors_io_out_23_Re),
    .io_out_23_Im(TwiddleFactors_io_out_23_Im),
    .io_out_24_Re(TwiddleFactors_io_out_24_Re),
    .io_out_24_Im(TwiddleFactors_io_out_24_Im),
    .io_out_25_Re(TwiddleFactors_io_out_25_Re),
    .io_out_25_Im(TwiddleFactors_io_out_25_Im),
    .io_out_26_Re(TwiddleFactors_io_out_26_Re),
    .io_out_26_Im(TwiddleFactors_io_out_26_Im),
    .io_out_27_Re(TwiddleFactors_io_out_27_Re),
    .io_out_27_Im(TwiddleFactors_io_out_27_Im),
    .io_out_28_Re(TwiddleFactors_io_out_28_Re),
    .io_out_28_Im(TwiddleFactors_io_out_28_Im),
    .io_out_29_Re(TwiddleFactors_io_out_29_Re),
    .io_out_29_Im(TwiddleFactors_io_out_29_Im),
    .io_out_30_Re(TwiddleFactors_io_out_30_Re),
    .io_out_30_Im(TwiddleFactors_io_out_30_Im),
    .io_out_31_Re(TwiddleFactors_io_out_31_Re),
    .io_out_31_Im(TwiddleFactors_io_out_31_Im)
  );
  TwiddleFactors_1 TwiddleFactors_1 ( // @[FFTDesigns.scala 3133:24]
    .clock(TwiddleFactors_1_clock),
    .reset(TwiddleFactors_1_reset),
    .io_in_0_Re(TwiddleFactors_1_io_in_0_Re),
    .io_in_0_Im(TwiddleFactors_1_io_in_0_Im),
    .io_in_1_Re(TwiddleFactors_1_io_in_1_Re),
    .io_in_1_Im(TwiddleFactors_1_io_in_1_Im),
    .io_in_2_Re(TwiddleFactors_1_io_in_2_Re),
    .io_in_2_Im(TwiddleFactors_1_io_in_2_Im),
    .io_in_3_Re(TwiddleFactors_1_io_in_3_Re),
    .io_in_3_Im(TwiddleFactors_1_io_in_3_Im),
    .io_in_4_Re(TwiddleFactors_1_io_in_4_Re),
    .io_in_4_Im(TwiddleFactors_1_io_in_4_Im),
    .io_in_5_Re(TwiddleFactors_1_io_in_5_Re),
    .io_in_5_Im(TwiddleFactors_1_io_in_5_Im),
    .io_in_6_Re(TwiddleFactors_1_io_in_6_Re),
    .io_in_6_Im(TwiddleFactors_1_io_in_6_Im),
    .io_in_7_Re(TwiddleFactors_1_io_in_7_Re),
    .io_in_7_Im(TwiddleFactors_1_io_in_7_Im),
    .io_in_8_Re(TwiddleFactors_1_io_in_8_Re),
    .io_in_8_Im(TwiddleFactors_1_io_in_8_Im),
    .io_in_9_Re(TwiddleFactors_1_io_in_9_Re),
    .io_in_9_Im(TwiddleFactors_1_io_in_9_Im),
    .io_in_10_Re(TwiddleFactors_1_io_in_10_Re),
    .io_in_10_Im(TwiddleFactors_1_io_in_10_Im),
    .io_in_11_Re(TwiddleFactors_1_io_in_11_Re),
    .io_in_11_Im(TwiddleFactors_1_io_in_11_Im),
    .io_in_12_Re(TwiddleFactors_1_io_in_12_Re),
    .io_in_12_Im(TwiddleFactors_1_io_in_12_Im),
    .io_in_13_Re(TwiddleFactors_1_io_in_13_Re),
    .io_in_13_Im(TwiddleFactors_1_io_in_13_Im),
    .io_in_14_Re(TwiddleFactors_1_io_in_14_Re),
    .io_in_14_Im(TwiddleFactors_1_io_in_14_Im),
    .io_in_15_Re(TwiddleFactors_1_io_in_15_Re),
    .io_in_15_Im(TwiddleFactors_1_io_in_15_Im),
    .io_in_16_Re(TwiddleFactors_1_io_in_16_Re),
    .io_in_16_Im(TwiddleFactors_1_io_in_16_Im),
    .io_in_17_Re(TwiddleFactors_1_io_in_17_Re),
    .io_in_17_Im(TwiddleFactors_1_io_in_17_Im),
    .io_in_18_Re(TwiddleFactors_1_io_in_18_Re),
    .io_in_18_Im(TwiddleFactors_1_io_in_18_Im),
    .io_in_19_Re(TwiddleFactors_1_io_in_19_Re),
    .io_in_19_Im(TwiddleFactors_1_io_in_19_Im),
    .io_in_20_Re(TwiddleFactors_1_io_in_20_Re),
    .io_in_20_Im(TwiddleFactors_1_io_in_20_Im),
    .io_in_21_Re(TwiddleFactors_1_io_in_21_Re),
    .io_in_21_Im(TwiddleFactors_1_io_in_21_Im),
    .io_in_22_Re(TwiddleFactors_1_io_in_22_Re),
    .io_in_22_Im(TwiddleFactors_1_io_in_22_Im),
    .io_in_23_Re(TwiddleFactors_1_io_in_23_Re),
    .io_in_23_Im(TwiddleFactors_1_io_in_23_Im),
    .io_in_24_Re(TwiddleFactors_1_io_in_24_Re),
    .io_in_24_Im(TwiddleFactors_1_io_in_24_Im),
    .io_in_25_Re(TwiddleFactors_1_io_in_25_Re),
    .io_in_25_Im(TwiddleFactors_1_io_in_25_Im),
    .io_in_26_Re(TwiddleFactors_1_io_in_26_Re),
    .io_in_26_Im(TwiddleFactors_1_io_in_26_Im),
    .io_in_27_Re(TwiddleFactors_1_io_in_27_Re),
    .io_in_27_Im(TwiddleFactors_1_io_in_27_Im),
    .io_in_28_Re(TwiddleFactors_1_io_in_28_Re),
    .io_in_28_Im(TwiddleFactors_1_io_in_28_Im),
    .io_in_29_Re(TwiddleFactors_1_io_in_29_Re),
    .io_in_29_Im(TwiddleFactors_1_io_in_29_Im),
    .io_in_30_Re(TwiddleFactors_1_io_in_30_Re),
    .io_in_30_Im(TwiddleFactors_1_io_in_30_Im),
    .io_in_31_Re(TwiddleFactors_1_io_in_31_Re),
    .io_in_31_Im(TwiddleFactors_1_io_in_31_Im),
    .io_out_0_Re(TwiddleFactors_1_io_out_0_Re),
    .io_out_0_Im(TwiddleFactors_1_io_out_0_Im),
    .io_out_1_Re(TwiddleFactors_1_io_out_1_Re),
    .io_out_1_Im(TwiddleFactors_1_io_out_1_Im),
    .io_out_2_Re(TwiddleFactors_1_io_out_2_Re),
    .io_out_2_Im(TwiddleFactors_1_io_out_2_Im),
    .io_out_3_Re(TwiddleFactors_1_io_out_3_Re),
    .io_out_3_Im(TwiddleFactors_1_io_out_3_Im),
    .io_out_4_Re(TwiddleFactors_1_io_out_4_Re),
    .io_out_4_Im(TwiddleFactors_1_io_out_4_Im),
    .io_out_5_Re(TwiddleFactors_1_io_out_5_Re),
    .io_out_5_Im(TwiddleFactors_1_io_out_5_Im),
    .io_out_6_Re(TwiddleFactors_1_io_out_6_Re),
    .io_out_6_Im(TwiddleFactors_1_io_out_6_Im),
    .io_out_7_Re(TwiddleFactors_1_io_out_7_Re),
    .io_out_7_Im(TwiddleFactors_1_io_out_7_Im),
    .io_out_8_Re(TwiddleFactors_1_io_out_8_Re),
    .io_out_8_Im(TwiddleFactors_1_io_out_8_Im),
    .io_out_9_Re(TwiddleFactors_1_io_out_9_Re),
    .io_out_9_Im(TwiddleFactors_1_io_out_9_Im),
    .io_out_10_Re(TwiddleFactors_1_io_out_10_Re),
    .io_out_10_Im(TwiddleFactors_1_io_out_10_Im),
    .io_out_11_Re(TwiddleFactors_1_io_out_11_Re),
    .io_out_11_Im(TwiddleFactors_1_io_out_11_Im),
    .io_out_12_Re(TwiddleFactors_1_io_out_12_Re),
    .io_out_12_Im(TwiddleFactors_1_io_out_12_Im),
    .io_out_13_Re(TwiddleFactors_1_io_out_13_Re),
    .io_out_13_Im(TwiddleFactors_1_io_out_13_Im),
    .io_out_14_Re(TwiddleFactors_1_io_out_14_Re),
    .io_out_14_Im(TwiddleFactors_1_io_out_14_Im),
    .io_out_15_Re(TwiddleFactors_1_io_out_15_Re),
    .io_out_15_Im(TwiddleFactors_1_io_out_15_Im),
    .io_out_16_Re(TwiddleFactors_1_io_out_16_Re),
    .io_out_16_Im(TwiddleFactors_1_io_out_16_Im),
    .io_out_17_Re(TwiddleFactors_1_io_out_17_Re),
    .io_out_17_Im(TwiddleFactors_1_io_out_17_Im),
    .io_out_18_Re(TwiddleFactors_1_io_out_18_Re),
    .io_out_18_Im(TwiddleFactors_1_io_out_18_Im),
    .io_out_19_Re(TwiddleFactors_1_io_out_19_Re),
    .io_out_19_Im(TwiddleFactors_1_io_out_19_Im),
    .io_out_20_Re(TwiddleFactors_1_io_out_20_Re),
    .io_out_20_Im(TwiddleFactors_1_io_out_20_Im),
    .io_out_21_Re(TwiddleFactors_1_io_out_21_Re),
    .io_out_21_Im(TwiddleFactors_1_io_out_21_Im),
    .io_out_22_Re(TwiddleFactors_1_io_out_22_Re),
    .io_out_22_Im(TwiddleFactors_1_io_out_22_Im),
    .io_out_23_Re(TwiddleFactors_1_io_out_23_Re),
    .io_out_23_Im(TwiddleFactors_1_io_out_23_Im),
    .io_out_24_Re(TwiddleFactors_1_io_out_24_Re),
    .io_out_24_Im(TwiddleFactors_1_io_out_24_Im),
    .io_out_25_Re(TwiddleFactors_1_io_out_25_Re),
    .io_out_25_Im(TwiddleFactors_1_io_out_25_Im),
    .io_out_26_Re(TwiddleFactors_1_io_out_26_Re),
    .io_out_26_Im(TwiddleFactors_1_io_out_26_Im),
    .io_out_27_Re(TwiddleFactors_1_io_out_27_Re),
    .io_out_27_Im(TwiddleFactors_1_io_out_27_Im),
    .io_out_28_Re(TwiddleFactors_1_io_out_28_Re),
    .io_out_28_Im(TwiddleFactors_1_io_out_28_Im),
    .io_out_29_Re(TwiddleFactors_1_io_out_29_Re),
    .io_out_29_Im(TwiddleFactors_1_io_out_29_Im),
    .io_out_30_Re(TwiddleFactors_1_io_out_30_Re),
    .io_out_30_Im(TwiddleFactors_1_io_out_30_Im),
    .io_out_31_Re(TwiddleFactors_1_io_out_31_Re),
    .io_out_31_Im(TwiddleFactors_1_io_out_31_Im)
  );
  TwiddleFactors_2 TwiddleFactors_2 ( // @[FFTDesigns.scala 3133:24]
    .clock(TwiddleFactors_2_clock),
    .reset(TwiddleFactors_2_reset),
    .io_in_0_Re(TwiddleFactors_2_io_in_0_Re),
    .io_in_0_Im(TwiddleFactors_2_io_in_0_Im),
    .io_in_1_Re(TwiddleFactors_2_io_in_1_Re),
    .io_in_1_Im(TwiddleFactors_2_io_in_1_Im),
    .io_in_2_Re(TwiddleFactors_2_io_in_2_Re),
    .io_in_2_Im(TwiddleFactors_2_io_in_2_Im),
    .io_in_3_Re(TwiddleFactors_2_io_in_3_Re),
    .io_in_3_Im(TwiddleFactors_2_io_in_3_Im),
    .io_in_4_Re(TwiddleFactors_2_io_in_4_Re),
    .io_in_4_Im(TwiddleFactors_2_io_in_4_Im),
    .io_in_5_Re(TwiddleFactors_2_io_in_5_Re),
    .io_in_5_Im(TwiddleFactors_2_io_in_5_Im),
    .io_in_6_Re(TwiddleFactors_2_io_in_6_Re),
    .io_in_6_Im(TwiddleFactors_2_io_in_6_Im),
    .io_in_7_Re(TwiddleFactors_2_io_in_7_Re),
    .io_in_7_Im(TwiddleFactors_2_io_in_7_Im),
    .io_in_8_Re(TwiddleFactors_2_io_in_8_Re),
    .io_in_8_Im(TwiddleFactors_2_io_in_8_Im),
    .io_in_9_Re(TwiddleFactors_2_io_in_9_Re),
    .io_in_9_Im(TwiddleFactors_2_io_in_9_Im),
    .io_in_10_Re(TwiddleFactors_2_io_in_10_Re),
    .io_in_10_Im(TwiddleFactors_2_io_in_10_Im),
    .io_in_11_Re(TwiddleFactors_2_io_in_11_Re),
    .io_in_11_Im(TwiddleFactors_2_io_in_11_Im),
    .io_in_12_Re(TwiddleFactors_2_io_in_12_Re),
    .io_in_12_Im(TwiddleFactors_2_io_in_12_Im),
    .io_in_13_Re(TwiddleFactors_2_io_in_13_Re),
    .io_in_13_Im(TwiddleFactors_2_io_in_13_Im),
    .io_in_14_Re(TwiddleFactors_2_io_in_14_Re),
    .io_in_14_Im(TwiddleFactors_2_io_in_14_Im),
    .io_in_15_Re(TwiddleFactors_2_io_in_15_Re),
    .io_in_15_Im(TwiddleFactors_2_io_in_15_Im),
    .io_in_16_Re(TwiddleFactors_2_io_in_16_Re),
    .io_in_16_Im(TwiddleFactors_2_io_in_16_Im),
    .io_in_17_Re(TwiddleFactors_2_io_in_17_Re),
    .io_in_17_Im(TwiddleFactors_2_io_in_17_Im),
    .io_in_18_Re(TwiddleFactors_2_io_in_18_Re),
    .io_in_18_Im(TwiddleFactors_2_io_in_18_Im),
    .io_in_19_Re(TwiddleFactors_2_io_in_19_Re),
    .io_in_19_Im(TwiddleFactors_2_io_in_19_Im),
    .io_in_20_Re(TwiddleFactors_2_io_in_20_Re),
    .io_in_20_Im(TwiddleFactors_2_io_in_20_Im),
    .io_in_21_Re(TwiddleFactors_2_io_in_21_Re),
    .io_in_21_Im(TwiddleFactors_2_io_in_21_Im),
    .io_in_22_Re(TwiddleFactors_2_io_in_22_Re),
    .io_in_22_Im(TwiddleFactors_2_io_in_22_Im),
    .io_in_23_Re(TwiddleFactors_2_io_in_23_Re),
    .io_in_23_Im(TwiddleFactors_2_io_in_23_Im),
    .io_in_24_Re(TwiddleFactors_2_io_in_24_Re),
    .io_in_24_Im(TwiddleFactors_2_io_in_24_Im),
    .io_in_25_Re(TwiddleFactors_2_io_in_25_Re),
    .io_in_25_Im(TwiddleFactors_2_io_in_25_Im),
    .io_in_26_Re(TwiddleFactors_2_io_in_26_Re),
    .io_in_26_Im(TwiddleFactors_2_io_in_26_Im),
    .io_in_27_Re(TwiddleFactors_2_io_in_27_Re),
    .io_in_27_Im(TwiddleFactors_2_io_in_27_Im),
    .io_in_28_Re(TwiddleFactors_2_io_in_28_Re),
    .io_in_28_Im(TwiddleFactors_2_io_in_28_Im),
    .io_in_29_Re(TwiddleFactors_2_io_in_29_Re),
    .io_in_29_Im(TwiddleFactors_2_io_in_29_Im),
    .io_in_30_Re(TwiddleFactors_2_io_in_30_Re),
    .io_in_30_Im(TwiddleFactors_2_io_in_30_Im),
    .io_in_31_Re(TwiddleFactors_2_io_in_31_Re),
    .io_in_31_Im(TwiddleFactors_2_io_in_31_Im),
    .io_out_0_Re(TwiddleFactors_2_io_out_0_Re),
    .io_out_0_Im(TwiddleFactors_2_io_out_0_Im),
    .io_out_1_Re(TwiddleFactors_2_io_out_1_Re),
    .io_out_1_Im(TwiddleFactors_2_io_out_1_Im),
    .io_out_2_Re(TwiddleFactors_2_io_out_2_Re),
    .io_out_2_Im(TwiddleFactors_2_io_out_2_Im),
    .io_out_3_Re(TwiddleFactors_2_io_out_3_Re),
    .io_out_3_Im(TwiddleFactors_2_io_out_3_Im),
    .io_out_4_Re(TwiddleFactors_2_io_out_4_Re),
    .io_out_4_Im(TwiddleFactors_2_io_out_4_Im),
    .io_out_5_Re(TwiddleFactors_2_io_out_5_Re),
    .io_out_5_Im(TwiddleFactors_2_io_out_5_Im),
    .io_out_6_Re(TwiddleFactors_2_io_out_6_Re),
    .io_out_6_Im(TwiddleFactors_2_io_out_6_Im),
    .io_out_7_Re(TwiddleFactors_2_io_out_7_Re),
    .io_out_7_Im(TwiddleFactors_2_io_out_7_Im),
    .io_out_8_Re(TwiddleFactors_2_io_out_8_Re),
    .io_out_8_Im(TwiddleFactors_2_io_out_8_Im),
    .io_out_9_Re(TwiddleFactors_2_io_out_9_Re),
    .io_out_9_Im(TwiddleFactors_2_io_out_9_Im),
    .io_out_10_Re(TwiddleFactors_2_io_out_10_Re),
    .io_out_10_Im(TwiddleFactors_2_io_out_10_Im),
    .io_out_11_Re(TwiddleFactors_2_io_out_11_Re),
    .io_out_11_Im(TwiddleFactors_2_io_out_11_Im),
    .io_out_12_Re(TwiddleFactors_2_io_out_12_Re),
    .io_out_12_Im(TwiddleFactors_2_io_out_12_Im),
    .io_out_13_Re(TwiddleFactors_2_io_out_13_Re),
    .io_out_13_Im(TwiddleFactors_2_io_out_13_Im),
    .io_out_14_Re(TwiddleFactors_2_io_out_14_Re),
    .io_out_14_Im(TwiddleFactors_2_io_out_14_Im),
    .io_out_15_Re(TwiddleFactors_2_io_out_15_Re),
    .io_out_15_Im(TwiddleFactors_2_io_out_15_Im),
    .io_out_16_Re(TwiddleFactors_2_io_out_16_Re),
    .io_out_16_Im(TwiddleFactors_2_io_out_16_Im),
    .io_out_17_Re(TwiddleFactors_2_io_out_17_Re),
    .io_out_17_Im(TwiddleFactors_2_io_out_17_Im),
    .io_out_18_Re(TwiddleFactors_2_io_out_18_Re),
    .io_out_18_Im(TwiddleFactors_2_io_out_18_Im),
    .io_out_19_Re(TwiddleFactors_2_io_out_19_Re),
    .io_out_19_Im(TwiddleFactors_2_io_out_19_Im),
    .io_out_20_Re(TwiddleFactors_2_io_out_20_Re),
    .io_out_20_Im(TwiddleFactors_2_io_out_20_Im),
    .io_out_21_Re(TwiddleFactors_2_io_out_21_Re),
    .io_out_21_Im(TwiddleFactors_2_io_out_21_Im),
    .io_out_22_Re(TwiddleFactors_2_io_out_22_Re),
    .io_out_22_Im(TwiddleFactors_2_io_out_22_Im),
    .io_out_23_Re(TwiddleFactors_2_io_out_23_Re),
    .io_out_23_Im(TwiddleFactors_2_io_out_23_Im),
    .io_out_24_Re(TwiddleFactors_2_io_out_24_Re),
    .io_out_24_Im(TwiddleFactors_2_io_out_24_Im),
    .io_out_25_Re(TwiddleFactors_2_io_out_25_Re),
    .io_out_25_Im(TwiddleFactors_2_io_out_25_Im),
    .io_out_26_Re(TwiddleFactors_2_io_out_26_Re),
    .io_out_26_Im(TwiddleFactors_2_io_out_26_Im),
    .io_out_27_Re(TwiddleFactors_2_io_out_27_Re),
    .io_out_27_Im(TwiddleFactors_2_io_out_27_Im),
    .io_out_28_Re(TwiddleFactors_2_io_out_28_Re),
    .io_out_28_Im(TwiddleFactors_2_io_out_28_Im),
    .io_out_29_Re(TwiddleFactors_2_io_out_29_Re),
    .io_out_29_Im(TwiddleFactors_2_io_out_29_Im),
    .io_out_30_Re(TwiddleFactors_2_io_out_30_Re),
    .io_out_30_Im(TwiddleFactors_2_io_out_30_Im),
    .io_out_31_Re(TwiddleFactors_2_io_out_31_Re),
    .io_out_31_Im(TwiddleFactors_2_io_out_31_Im)
  );
  TwiddleFactors_3 TwiddleFactors_3 ( // @[FFTDesigns.scala 3133:24]
    .clock(TwiddleFactors_3_clock),
    .reset(TwiddleFactors_3_reset),
    .io_in_0_Re(TwiddleFactors_3_io_in_0_Re),
    .io_in_0_Im(TwiddleFactors_3_io_in_0_Im),
    .io_in_1_Re(TwiddleFactors_3_io_in_1_Re),
    .io_in_1_Im(TwiddleFactors_3_io_in_1_Im),
    .io_in_2_Re(TwiddleFactors_3_io_in_2_Re),
    .io_in_2_Im(TwiddleFactors_3_io_in_2_Im),
    .io_in_3_Re(TwiddleFactors_3_io_in_3_Re),
    .io_in_3_Im(TwiddleFactors_3_io_in_3_Im),
    .io_in_4_Re(TwiddleFactors_3_io_in_4_Re),
    .io_in_4_Im(TwiddleFactors_3_io_in_4_Im),
    .io_in_5_Re(TwiddleFactors_3_io_in_5_Re),
    .io_in_5_Im(TwiddleFactors_3_io_in_5_Im),
    .io_in_6_Re(TwiddleFactors_3_io_in_6_Re),
    .io_in_6_Im(TwiddleFactors_3_io_in_6_Im),
    .io_in_7_Re(TwiddleFactors_3_io_in_7_Re),
    .io_in_7_Im(TwiddleFactors_3_io_in_7_Im),
    .io_in_8_Re(TwiddleFactors_3_io_in_8_Re),
    .io_in_8_Im(TwiddleFactors_3_io_in_8_Im),
    .io_in_9_Re(TwiddleFactors_3_io_in_9_Re),
    .io_in_9_Im(TwiddleFactors_3_io_in_9_Im),
    .io_in_10_Re(TwiddleFactors_3_io_in_10_Re),
    .io_in_10_Im(TwiddleFactors_3_io_in_10_Im),
    .io_in_11_Re(TwiddleFactors_3_io_in_11_Re),
    .io_in_11_Im(TwiddleFactors_3_io_in_11_Im),
    .io_in_12_Re(TwiddleFactors_3_io_in_12_Re),
    .io_in_12_Im(TwiddleFactors_3_io_in_12_Im),
    .io_in_13_Re(TwiddleFactors_3_io_in_13_Re),
    .io_in_13_Im(TwiddleFactors_3_io_in_13_Im),
    .io_in_14_Re(TwiddleFactors_3_io_in_14_Re),
    .io_in_14_Im(TwiddleFactors_3_io_in_14_Im),
    .io_in_15_Re(TwiddleFactors_3_io_in_15_Re),
    .io_in_15_Im(TwiddleFactors_3_io_in_15_Im),
    .io_in_16_Re(TwiddleFactors_3_io_in_16_Re),
    .io_in_16_Im(TwiddleFactors_3_io_in_16_Im),
    .io_in_17_Re(TwiddleFactors_3_io_in_17_Re),
    .io_in_17_Im(TwiddleFactors_3_io_in_17_Im),
    .io_in_18_Re(TwiddleFactors_3_io_in_18_Re),
    .io_in_18_Im(TwiddleFactors_3_io_in_18_Im),
    .io_in_19_Re(TwiddleFactors_3_io_in_19_Re),
    .io_in_19_Im(TwiddleFactors_3_io_in_19_Im),
    .io_in_20_Re(TwiddleFactors_3_io_in_20_Re),
    .io_in_20_Im(TwiddleFactors_3_io_in_20_Im),
    .io_in_21_Re(TwiddleFactors_3_io_in_21_Re),
    .io_in_21_Im(TwiddleFactors_3_io_in_21_Im),
    .io_in_22_Re(TwiddleFactors_3_io_in_22_Re),
    .io_in_22_Im(TwiddleFactors_3_io_in_22_Im),
    .io_in_23_Re(TwiddleFactors_3_io_in_23_Re),
    .io_in_23_Im(TwiddleFactors_3_io_in_23_Im),
    .io_in_24_Re(TwiddleFactors_3_io_in_24_Re),
    .io_in_24_Im(TwiddleFactors_3_io_in_24_Im),
    .io_in_25_Re(TwiddleFactors_3_io_in_25_Re),
    .io_in_25_Im(TwiddleFactors_3_io_in_25_Im),
    .io_in_26_Re(TwiddleFactors_3_io_in_26_Re),
    .io_in_26_Im(TwiddleFactors_3_io_in_26_Im),
    .io_in_27_Re(TwiddleFactors_3_io_in_27_Re),
    .io_in_27_Im(TwiddleFactors_3_io_in_27_Im),
    .io_in_28_Re(TwiddleFactors_3_io_in_28_Re),
    .io_in_28_Im(TwiddleFactors_3_io_in_28_Im),
    .io_in_29_Re(TwiddleFactors_3_io_in_29_Re),
    .io_in_29_Im(TwiddleFactors_3_io_in_29_Im),
    .io_in_30_Re(TwiddleFactors_3_io_in_30_Re),
    .io_in_30_Im(TwiddleFactors_3_io_in_30_Im),
    .io_in_31_Re(TwiddleFactors_3_io_in_31_Re),
    .io_in_31_Im(TwiddleFactors_3_io_in_31_Im),
    .io_out_0_Re(TwiddleFactors_3_io_out_0_Re),
    .io_out_0_Im(TwiddleFactors_3_io_out_0_Im),
    .io_out_1_Re(TwiddleFactors_3_io_out_1_Re),
    .io_out_1_Im(TwiddleFactors_3_io_out_1_Im),
    .io_out_2_Re(TwiddleFactors_3_io_out_2_Re),
    .io_out_2_Im(TwiddleFactors_3_io_out_2_Im),
    .io_out_3_Re(TwiddleFactors_3_io_out_3_Re),
    .io_out_3_Im(TwiddleFactors_3_io_out_3_Im),
    .io_out_4_Re(TwiddleFactors_3_io_out_4_Re),
    .io_out_4_Im(TwiddleFactors_3_io_out_4_Im),
    .io_out_5_Re(TwiddleFactors_3_io_out_5_Re),
    .io_out_5_Im(TwiddleFactors_3_io_out_5_Im),
    .io_out_6_Re(TwiddleFactors_3_io_out_6_Re),
    .io_out_6_Im(TwiddleFactors_3_io_out_6_Im),
    .io_out_7_Re(TwiddleFactors_3_io_out_7_Re),
    .io_out_7_Im(TwiddleFactors_3_io_out_7_Im),
    .io_out_8_Re(TwiddleFactors_3_io_out_8_Re),
    .io_out_8_Im(TwiddleFactors_3_io_out_8_Im),
    .io_out_9_Re(TwiddleFactors_3_io_out_9_Re),
    .io_out_9_Im(TwiddleFactors_3_io_out_9_Im),
    .io_out_10_Re(TwiddleFactors_3_io_out_10_Re),
    .io_out_10_Im(TwiddleFactors_3_io_out_10_Im),
    .io_out_11_Re(TwiddleFactors_3_io_out_11_Re),
    .io_out_11_Im(TwiddleFactors_3_io_out_11_Im),
    .io_out_12_Re(TwiddleFactors_3_io_out_12_Re),
    .io_out_12_Im(TwiddleFactors_3_io_out_12_Im),
    .io_out_13_Re(TwiddleFactors_3_io_out_13_Re),
    .io_out_13_Im(TwiddleFactors_3_io_out_13_Im),
    .io_out_14_Re(TwiddleFactors_3_io_out_14_Re),
    .io_out_14_Im(TwiddleFactors_3_io_out_14_Im),
    .io_out_15_Re(TwiddleFactors_3_io_out_15_Re),
    .io_out_15_Im(TwiddleFactors_3_io_out_15_Im),
    .io_out_16_Re(TwiddleFactors_3_io_out_16_Re),
    .io_out_16_Im(TwiddleFactors_3_io_out_16_Im),
    .io_out_17_Re(TwiddleFactors_3_io_out_17_Re),
    .io_out_17_Im(TwiddleFactors_3_io_out_17_Im),
    .io_out_18_Re(TwiddleFactors_3_io_out_18_Re),
    .io_out_18_Im(TwiddleFactors_3_io_out_18_Im),
    .io_out_19_Re(TwiddleFactors_3_io_out_19_Re),
    .io_out_19_Im(TwiddleFactors_3_io_out_19_Im),
    .io_out_20_Re(TwiddleFactors_3_io_out_20_Re),
    .io_out_20_Im(TwiddleFactors_3_io_out_20_Im),
    .io_out_21_Re(TwiddleFactors_3_io_out_21_Re),
    .io_out_21_Im(TwiddleFactors_3_io_out_21_Im),
    .io_out_22_Re(TwiddleFactors_3_io_out_22_Re),
    .io_out_22_Im(TwiddleFactors_3_io_out_22_Im),
    .io_out_23_Re(TwiddleFactors_3_io_out_23_Re),
    .io_out_23_Im(TwiddleFactors_3_io_out_23_Im),
    .io_out_24_Re(TwiddleFactors_3_io_out_24_Re),
    .io_out_24_Im(TwiddleFactors_3_io_out_24_Im),
    .io_out_25_Re(TwiddleFactors_3_io_out_25_Re),
    .io_out_25_Im(TwiddleFactors_3_io_out_25_Im),
    .io_out_26_Re(TwiddleFactors_3_io_out_26_Re),
    .io_out_26_Im(TwiddleFactors_3_io_out_26_Im),
    .io_out_27_Re(TwiddleFactors_3_io_out_27_Re),
    .io_out_27_Im(TwiddleFactors_3_io_out_27_Im),
    .io_out_28_Re(TwiddleFactors_3_io_out_28_Re),
    .io_out_28_Im(TwiddleFactors_3_io_out_28_Im),
    .io_out_29_Re(TwiddleFactors_3_io_out_29_Re),
    .io_out_29_Im(TwiddleFactors_3_io_out_29_Im),
    .io_out_30_Re(TwiddleFactors_3_io_out_30_Re),
    .io_out_30_Im(TwiddleFactors_3_io_out_30_Im),
    .io_out_31_Re(TwiddleFactors_3_io_out_31_Re),
    .io_out_31_Im(TwiddleFactors_3_io_out_31_Im)
  );
  assign io_out_0_Re = PermutationsBasic_5_io_out_0_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_0_Im = PermutationsBasic_5_io_out_0_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_1_Re = PermutationsBasic_5_io_out_1_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_1_Im = PermutationsBasic_5_io_out_1_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_2_Re = PermutationsBasic_5_io_out_2_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_2_Im = PermutationsBasic_5_io_out_2_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_3_Re = PermutationsBasic_5_io_out_3_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_3_Im = PermutationsBasic_5_io_out_3_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_4_Re = PermutationsBasic_5_io_out_4_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_4_Im = PermutationsBasic_5_io_out_4_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_5_Re = PermutationsBasic_5_io_out_5_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_5_Im = PermutationsBasic_5_io_out_5_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_6_Re = PermutationsBasic_5_io_out_6_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_6_Im = PermutationsBasic_5_io_out_6_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_7_Re = PermutationsBasic_5_io_out_7_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_7_Im = PermutationsBasic_5_io_out_7_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_8_Re = PermutationsBasic_5_io_out_8_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_8_Im = PermutationsBasic_5_io_out_8_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_9_Re = PermutationsBasic_5_io_out_9_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_9_Im = PermutationsBasic_5_io_out_9_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_10_Re = PermutationsBasic_5_io_out_10_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_10_Im = PermutationsBasic_5_io_out_10_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_11_Re = PermutationsBasic_5_io_out_11_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_11_Im = PermutationsBasic_5_io_out_11_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_12_Re = PermutationsBasic_5_io_out_12_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_12_Im = PermutationsBasic_5_io_out_12_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_13_Re = PermutationsBasic_5_io_out_13_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_13_Im = PermutationsBasic_5_io_out_13_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_14_Re = PermutationsBasic_5_io_out_14_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_14_Im = PermutationsBasic_5_io_out_14_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_15_Re = PermutationsBasic_5_io_out_15_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_15_Im = PermutationsBasic_5_io_out_15_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_16_Re = PermutationsBasic_5_io_out_16_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_16_Im = PermutationsBasic_5_io_out_16_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_17_Re = PermutationsBasic_5_io_out_17_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_17_Im = PermutationsBasic_5_io_out_17_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_18_Re = PermutationsBasic_5_io_out_18_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_18_Im = PermutationsBasic_5_io_out_18_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_19_Re = PermutationsBasic_5_io_out_19_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_19_Im = PermutationsBasic_5_io_out_19_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_20_Re = PermutationsBasic_5_io_out_20_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_20_Im = PermutationsBasic_5_io_out_20_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_21_Re = PermutationsBasic_5_io_out_21_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_21_Im = PermutationsBasic_5_io_out_21_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_22_Re = PermutationsBasic_5_io_out_22_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_22_Im = PermutationsBasic_5_io_out_22_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_23_Re = PermutationsBasic_5_io_out_23_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_23_Im = PermutationsBasic_5_io_out_23_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_24_Re = PermutationsBasic_5_io_out_24_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_24_Im = PermutationsBasic_5_io_out_24_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_25_Re = PermutationsBasic_5_io_out_25_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_25_Im = PermutationsBasic_5_io_out_25_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_26_Re = PermutationsBasic_5_io_out_26_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_26_Im = PermutationsBasic_5_io_out_26_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_27_Re = PermutationsBasic_5_io_out_27_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_27_Im = PermutationsBasic_5_io_out_27_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_28_Re = PermutationsBasic_5_io_out_28_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_28_Im = PermutationsBasic_5_io_out_28_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_29_Re = PermutationsBasic_5_io_out_29_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_29_Im = PermutationsBasic_5_io_out_29_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_30_Re = PermutationsBasic_5_io_out_30_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_30_Im = PermutationsBasic_5_io_out_30_Im; // @[FFTDesigns.scala 3159:12]
  assign io_out_31_Re = PermutationsBasic_5_io_out_31_Re; // @[FFTDesigns.scala 3159:12]
  assign io_out_31_Im = PermutationsBasic_5_io_out_31_Im; // @[FFTDesigns.scala 3159:12]
  assign DFT_r_v2_clock = clock;
  assign DFT_r_v2_reset = reset;
  assign DFT_r_v2_io_in_0_Re = PermutationsBasic_io_out_0_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_io_in_0_Im = PermutationsBasic_io_out_0_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_io_in_1_Re = PermutationsBasic_io_out_1_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_io_in_1_Im = PermutationsBasic_io_out_1_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_1_clock = clock;
  assign DFT_r_v2_1_reset = reset;
  assign DFT_r_v2_1_io_in_0_Re = PermutationsBasic_io_out_2_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_1_io_in_0_Im = PermutationsBasic_io_out_2_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_1_io_in_1_Re = PermutationsBasic_io_out_3_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_1_io_in_1_Im = PermutationsBasic_io_out_3_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_2_clock = clock;
  assign DFT_r_v2_2_reset = reset;
  assign DFT_r_v2_2_io_in_0_Re = PermutationsBasic_io_out_4_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_2_io_in_0_Im = PermutationsBasic_io_out_4_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_2_io_in_1_Re = PermutationsBasic_io_out_5_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_2_io_in_1_Im = PermutationsBasic_io_out_5_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_3_clock = clock;
  assign DFT_r_v2_3_reset = reset;
  assign DFT_r_v2_3_io_in_0_Re = PermutationsBasic_io_out_6_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_3_io_in_0_Im = PermutationsBasic_io_out_6_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_3_io_in_1_Re = PermutationsBasic_io_out_7_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_3_io_in_1_Im = PermutationsBasic_io_out_7_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_4_clock = clock;
  assign DFT_r_v2_4_reset = reset;
  assign DFT_r_v2_4_io_in_0_Re = PermutationsBasic_io_out_8_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_4_io_in_0_Im = PermutationsBasic_io_out_8_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_4_io_in_1_Re = PermutationsBasic_io_out_9_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_4_io_in_1_Im = PermutationsBasic_io_out_9_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_5_clock = clock;
  assign DFT_r_v2_5_reset = reset;
  assign DFT_r_v2_5_io_in_0_Re = PermutationsBasic_io_out_10_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_5_io_in_0_Im = PermutationsBasic_io_out_10_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_5_io_in_1_Re = PermutationsBasic_io_out_11_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_5_io_in_1_Im = PermutationsBasic_io_out_11_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_6_clock = clock;
  assign DFT_r_v2_6_reset = reset;
  assign DFT_r_v2_6_io_in_0_Re = PermutationsBasic_io_out_12_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_6_io_in_0_Im = PermutationsBasic_io_out_12_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_6_io_in_1_Re = PermutationsBasic_io_out_13_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_6_io_in_1_Im = PermutationsBasic_io_out_13_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_7_clock = clock;
  assign DFT_r_v2_7_reset = reset;
  assign DFT_r_v2_7_io_in_0_Re = PermutationsBasic_io_out_14_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_7_io_in_0_Im = PermutationsBasic_io_out_14_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_7_io_in_1_Re = PermutationsBasic_io_out_15_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_7_io_in_1_Im = PermutationsBasic_io_out_15_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_8_clock = clock;
  assign DFT_r_v2_8_reset = reset;
  assign DFT_r_v2_8_io_in_0_Re = PermutationsBasic_io_out_16_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_8_io_in_0_Im = PermutationsBasic_io_out_16_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_8_io_in_1_Re = PermutationsBasic_io_out_17_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_8_io_in_1_Im = PermutationsBasic_io_out_17_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_9_clock = clock;
  assign DFT_r_v2_9_reset = reset;
  assign DFT_r_v2_9_io_in_0_Re = PermutationsBasic_io_out_18_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_9_io_in_0_Im = PermutationsBasic_io_out_18_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_9_io_in_1_Re = PermutationsBasic_io_out_19_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_9_io_in_1_Im = PermutationsBasic_io_out_19_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_10_clock = clock;
  assign DFT_r_v2_10_reset = reset;
  assign DFT_r_v2_10_io_in_0_Re = PermutationsBasic_io_out_20_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_10_io_in_0_Im = PermutationsBasic_io_out_20_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_10_io_in_1_Re = PermutationsBasic_io_out_21_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_10_io_in_1_Im = PermutationsBasic_io_out_21_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_11_clock = clock;
  assign DFT_r_v2_11_reset = reset;
  assign DFT_r_v2_11_io_in_0_Re = PermutationsBasic_io_out_22_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_11_io_in_0_Im = PermutationsBasic_io_out_22_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_11_io_in_1_Re = PermutationsBasic_io_out_23_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_11_io_in_1_Im = PermutationsBasic_io_out_23_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_12_clock = clock;
  assign DFT_r_v2_12_reset = reset;
  assign DFT_r_v2_12_io_in_0_Re = PermutationsBasic_io_out_24_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_12_io_in_0_Im = PermutationsBasic_io_out_24_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_12_io_in_1_Re = PermutationsBasic_io_out_25_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_12_io_in_1_Im = PermutationsBasic_io_out_25_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_13_clock = clock;
  assign DFT_r_v2_13_reset = reset;
  assign DFT_r_v2_13_io_in_0_Re = PermutationsBasic_io_out_26_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_13_io_in_0_Im = PermutationsBasic_io_out_26_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_13_io_in_1_Re = PermutationsBasic_io_out_27_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_13_io_in_1_Im = PermutationsBasic_io_out_27_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_14_clock = clock;
  assign DFT_r_v2_14_reset = reset;
  assign DFT_r_v2_14_io_in_0_Re = PermutationsBasic_io_out_28_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_14_io_in_0_Im = PermutationsBasic_io_out_28_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_14_io_in_1_Re = PermutationsBasic_io_out_29_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_14_io_in_1_Im = PermutationsBasic_io_out_29_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_15_clock = clock;
  assign DFT_r_v2_15_reset = reset;
  assign DFT_r_v2_15_io_in_0_Re = PermutationsBasic_io_out_30_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_15_io_in_0_Im = PermutationsBasic_io_out_30_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_15_io_in_1_Re = PermutationsBasic_io_out_31_Re; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_15_io_in_1_Im = PermutationsBasic_io_out_31_Im; // @[FFTDesigns.scala 3145:39]
  assign DFT_r_v2_16_clock = clock;
  assign DFT_r_v2_16_reset = reset;
  assign DFT_r_v2_16_io_in_0_Re = TwiddleFactors_io_out_0_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_16_io_in_0_Im = TwiddleFactors_io_out_0_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_16_io_in_1_Re = TwiddleFactors_io_out_1_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_16_io_in_1_Im = TwiddleFactors_io_out_1_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_17_clock = clock;
  assign DFT_r_v2_17_reset = reset;
  assign DFT_r_v2_17_io_in_0_Re = TwiddleFactors_io_out_2_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_17_io_in_0_Im = TwiddleFactors_io_out_2_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_17_io_in_1_Re = TwiddleFactors_io_out_3_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_17_io_in_1_Im = TwiddleFactors_io_out_3_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_18_clock = clock;
  assign DFT_r_v2_18_reset = reset;
  assign DFT_r_v2_18_io_in_0_Re = TwiddleFactors_io_out_4_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_18_io_in_0_Im = TwiddleFactors_io_out_4_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_18_io_in_1_Re = TwiddleFactors_io_out_5_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_18_io_in_1_Im = TwiddleFactors_io_out_5_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_19_clock = clock;
  assign DFT_r_v2_19_reset = reset;
  assign DFT_r_v2_19_io_in_0_Re = TwiddleFactors_io_out_6_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_19_io_in_0_Im = TwiddleFactors_io_out_6_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_19_io_in_1_Re = TwiddleFactors_io_out_7_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_19_io_in_1_Im = TwiddleFactors_io_out_7_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_20_clock = clock;
  assign DFT_r_v2_20_reset = reset;
  assign DFT_r_v2_20_io_in_0_Re = TwiddleFactors_io_out_8_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_20_io_in_0_Im = TwiddleFactors_io_out_8_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_20_io_in_1_Re = TwiddleFactors_io_out_9_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_20_io_in_1_Im = TwiddleFactors_io_out_9_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_21_clock = clock;
  assign DFT_r_v2_21_reset = reset;
  assign DFT_r_v2_21_io_in_0_Re = TwiddleFactors_io_out_10_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_21_io_in_0_Im = TwiddleFactors_io_out_10_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_21_io_in_1_Re = TwiddleFactors_io_out_11_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_21_io_in_1_Im = TwiddleFactors_io_out_11_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_22_clock = clock;
  assign DFT_r_v2_22_reset = reset;
  assign DFT_r_v2_22_io_in_0_Re = TwiddleFactors_io_out_12_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_22_io_in_0_Im = TwiddleFactors_io_out_12_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_22_io_in_1_Re = TwiddleFactors_io_out_13_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_22_io_in_1_Im = TwiddleFactors_io_out_13_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_23_clock = clock;
  assign DFT_r_v2_23_reset = reset;
  assign DFT_r_v2_23_io_in_0_Re = TwiddleFactors_io_out_14_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_23_io_in_0_Im = TwiddleFactors_io_out_14_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_23_io_in_1_Re = TwiddleFactors_io_out_15_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_23_io_in_1_Im = TwiddleFactors_io_out_15_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_24_clock = clock;
  assign DFT_r_v2_24_reset = reset;
  assign DFT_r_v2_24_io_in_0_Re = TwiddleFactors_io_out_16_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_24_io_in_0_Im = TwiddleFactors_io_out_16_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_24_io_in_1_Re = TwiddleFactors_io_out_17_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_24_io_in_1_Im = TwiddleFactors_io_out_17_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_25_clock = clock;
  assign DFT_r_v2_25_reset = reset;
  assign DFT_r_v2_25_io_in_0_Re = TwiddleFactors_io_out_18_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_25_io_in_0_Im = TwiddleFactors_io_out_18_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_25_io_in_1_Re = TwiddleFactors_io_out_19_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_25_io_in_1_Im = TwiddleFactors_io_out_19_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_26_clock = clock;
  assign DFT_r_v2_26_reset = reset;
  assign DFT_r_v2_26_io_in_0_Re = TwiddleFactors_io_out_20_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_26_io_in_0_Im = TwiddleFactors_io_out_20_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_26_io_in_1_Re = TwiddleFactors_io_out_21_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_26_io_in_1_Im = TwiddleFactors_io_out_21_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_27_clock = clock;
  assign DFT_r_v2_27_reset = reset;
  assign DFT_r_v2_27_io_in_0_Re = TwiddleFactors_io_out_22_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_27_io_in_0_Im = TwiddleFactors_io_out_22_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_27_io_in_1_Re = TwiddleFactors_io_out_23_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_27_io_in_1_Im = TwiddleFactors_io_out_23_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_28_clock = clock;
  assign DFT_r_v2_28_reset = reset;
  assign DFT_r_v2_28_io_in_0_Re = TwiddleFactors_io_out_24_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_28_io_in_0_Im = TwiddleFactors_io_out_24_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_28_io_in_1_Re = TwiddleFactors_io_out_25_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_28_io_in_1_Im = TwiddleFactors_io_out_25_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_29_clock = clock;
  assign DFT_r_v2_29_reset = reset;
  assign DFT_r_v2_29_io_in_0_Re = TwiddleFactors_io_out_26_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_29_io_in_0_Im = TwiddleFactors_io_out_26_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_29_io_in_1_Re = TwiddleFactors_io_out_27_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_29_io_in_1_Im = TwiddleFactors_io_out_27_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_30_clock = clock;
  assign DFT_r_v2_30_reset = reset;
  assign DFT_r_v2_30_io_in_0_Re = TwiddleFactors_io_out_28_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_30_io_in_0_Im = TwiddleFactors_io_out_28_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_30_io_in_1_Re = TwiddleFactors_io_out_29_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_30_io_in_1_Im = TwiddleFactors_io_out_29_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_31_clock = clock;
  assign DFT_r_v2_31_reset = reset;
  assign DFT_r_v2_31_io_in_0_Re = TwiddleFactors_io_out_30_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_31_io_in_0_Im = TwiddleFactors_io_out_30_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_31_io_in_1_Re = TwiddleFactors_io_out_31_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_31_io_in_1_Im = TwiddleFactors_io_out_31_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_32_clock = clock;
  assign DFT_r_v2_32_reset = reset;
  assign DFT_r_v2_32_io_in_0_Re = TwiddleFactors_1_io_out_0_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_32_io_in_0_Im = TwiddleFactors_1_io_out_0_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_32_io_in_1_Re = TwiddleFactors_1_io_out_1_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_32_io_in_1_Im = TwiddleFactors_1_io_out_1_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_33_clock = clock;
  assign DFT_r_v2_33_reset = reset;
  assign DFT_r_v2_33_io_in_0_Re = TwiddleFactors_1_io_out_2_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_33_io_in_0_Im = TwiddleFactors_1_io_out_2_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_33_io_in_1_Re = TwiddleFactors_1_io_out_3_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_33_io_in_1_Im = TwiddleFactors_1_io_out_3_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_34_clock = clock;
  assign DFT_r_v2_34_reset = reset;
  assign DFT_r_v2_34_io_in_0_Re = TwiddleFactors_1_io_out_4_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_34_io_in_0_Im = TwiddleFactors_1_io_out_4_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_34_io_in_1_Re = TwiddleFactors_1_io_out_5_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_34_io_in_1_Im = TwiddleFactors_1_io_out_5_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_35_clock = clock;
  assign DFT_r_v2_35_reset = reset;
  assign DFT_r_v2_35_io_in_0_Re = TwiddleFactors_1_io_out_6_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_35_io_in_0_Im = TwiddleFactors_1_io_out_6_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_35_io_in_1_Re = TwiddleFactors_1_io_out_7_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_35_io_in_1_Im = TwiddleFactors_1_io_out_7_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_36_clock = clock;
  assign DFT_r_v2_36_reset = reset;
  assign DFT_r_v2_36_io_in_0_Re = TwiddleFactors_1_io_out_8_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_36_io_in_0_Im = TwiddleFactors_1_io_out_8_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_36_io_in_1_Re = TwiddleFactors_1_io_out_9_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_36_io_in_1_Im = TwiddleFactors_1_io_out_9_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_37_clock = clock;
  assign DFT_r_v2_37_reset = reset;
  assign DFT_r_v2_37_io_in_0_Re = TwiddleFactors_1_io_out_10_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_37_io_in_0_Im = TwiddleFactors_1_io_out_10_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_37_io_in_1_Re = TwiddleFactors_1_io_out_11_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_37_io_in_1_Im = TwiddleFactors_1_io_out_11_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_38_clock = clock;
  assign DFT_r_v2_38_reset = reset;
  assign DFT_r_v2_38_io_in_0_Re = TwiddleFactors_1_io_out_12_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_38_io_in_0_Im = TwiddleFactors_1_io_out_12_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_38_io_in_1_Re = TwiddleFactors_1_io_out_13_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_38_io_in_1_Im = TwiddleFactors_1_io_out_13_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_39_clock = clock;
  assign DFT_r_v2_39_reset = reset;
  assign DFT_r_v2_39_io_in_0_Re = TwiddleFactors_1_io_out_14_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_39_io_in_0_Im = TwiddleFactors_1_io_out_14_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_39_io_in_1_Re = TwiddleFactors_1_io_out_15_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_39_io_in_1_Im = TwiddleFactors_1_io_out_15_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_40_clock = clock;
  assign DFT_r_v2_40_reset = reset;
  assign DFT_r_v2_40_io_in_0_Re = TwiddleFactors_1_io_out_16_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_40_io_in_0_Im = TwiddleFactors_1_io_out_16_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_40_io_in_1_Re = TwiddleFactors_1_io_out_17_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_40_io_in_1_Im = TwiddleFactors_1_io_out_17_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_41_clock = clock;
  assign DFT_r_v2_41_reset = reset;
  assign DFT_r_v2_41_io_in_0_Re = TwiddleFactors_1_io_out_18_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_41_io_in_0_Im = TwiddleFactors_1_io_out_18_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_41_io_in_1_Re = TwiddleFactors_1_io_out_19_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_41_io_in_1_Im = TwiddleFactors_1_io_out_19_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_42_clock = clock;
  assign DFT_r_v2_42_reset = reset;
  assign DFT_r_v2_42_io_in_0_Re = TwiddleFactors_1_io_out_20_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_42_io_in_0_Im = TwiddleFactors_1_io_out_20_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_42_io_in_1_Re = TwiddleFactors_1_io_out_21_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_42_io_in_1_Im = TwiddleFactors_1_io_out_21_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_43_clock = clock;
  assign DFT_r_v2_43_reset = reset;
  assign DFT_r_v2_43_io_in_0_Re = TwiddleFactors_1_io_out_22_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_43_io_in_0_Im = TwiddleFactors_1_io_out_22_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_43_io_in_1_Re = TwiddleFactors_1_io_out_23_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_43_io_in_1_Im = TwiddleFactors_1_io_out_23_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_44_clock = clock;
  assign DFT_r_v2_44_reset = reset;
  assign DFT_r_v2_44_io_in_0_Re = TwiddleFactors_1_io_out_24_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_44_io_in_0_Im = TwiddleFactors_1_io_out_24_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_44_io_in_1_Re = TwiddleFactors_1_io_out_25_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_44_io_in_1_Im = TwiddleFactors_1_io_out_25_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_45_clock = clock;
  assign DFT_r_v2_45_reset = reset;
  assign DFT_r_v2_45_io_in_0_Re = TwiddleFactors_1_io_out_26_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_45_io_in_0_Im = TwiddleFactors_1_io_out_26_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_45_io_in_1_Re = TwiddleFactors_1_io_out_27_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_45_io_in_1_Im = TwiddleFactors_1_io_out_27_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_46_clock = clock;
  assign DFT_r_v2_46_reset = reset;
  assign DFT_r_v2_46_io_in_0_Re = TwiddleFactors_1_io_out_28_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_46_io_in_0_Im = TwiddleFactors_1_io_out_28_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_46_io_in_1_Re = TwiddleFactors_1_io_out_29_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_46_io_in_1_Im = TwiddleFactors_1_io_out_29_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_47_clock = clock;
  assign DFT_r_v2_47_reset = reset;
  assign DFT_r_v2_47_io_in_0_Re = TwiddleFactors_1_io_out_30_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_47_io_in_0_Im = TwiddleFactors_1_io_out_30_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_47_io_in_1_Re = TwiddleFactors_1_io_out_31_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_47_io_in_1_Im = TwiddleFactors_1_io_out_31_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_48_clock = clock;
  assign DFT_r_v2_48_reset = reset;
  assign DFT_r_v2_48_io_in_0_Re = TwiddleFactors_2_io_out_0_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_48_io_in_0_Im = TwiddleFactors_2_io_out_0_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_48_io_in_1_Re = TwiddleFactors_2_io_out_1_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_48_io_in_1_Im = TwiddleFactors_2_io_out_1_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_49_clock = clock;
  assign DFT_r_v2_49_reset = reset;
  assign DFT_r_v2_49_io_in_0_Re = TwiddleFactors_2_io_out_2_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_49_io_in_0_Im = TwiddleFactors_2_io_out_2_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_49_io_in_1_Re = TwiddleFactors_2_io_out_3_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_49_io_in_1_Im = TwiddleFactors_2_io_out_3_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_50_clock = clock;
  assign DFT_r_v2_50_reset = reset;
  assign DFT_r_v2_50_io_in_0_Re = TwiddleFactors_2_io_out_4_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_50_io_in_0_Im = TwiddleFactors_2_io_out_4_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_50_io_in_1_Re = TwiddleFactors_2_io_out_5_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_50_io_in_1_Im = TwiddleFactors_2_io_out_5_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_51_clock = clock;
  assign DFT_r_v2_51_reset = reset;
  assign DFT_r_v2_51_io_in_0_Re = TwiddleFactors_2_io_out_6_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_51_io_in_0_Im = TwiddleFactors_2_io_out_6_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_51_io_in_1_Re = TwiddleFactors_2_io_out_7_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_51_io_in_1_Im = TwiddleFactors_2_io_out_7_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_52_clock = clock;
  assign DFT_r_v2_52_reset = reset;
  assign DFT_r_v2_52_io_in_0_Re = TwiddleFactors_2_io_out_8_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_52_io_in_0_Im = TwiddleFactors_2_io_out_8_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_52_io_in_1_Re = TwiddleFactors_2_io_out_9_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_52_io_in_1_Im = TwiddleFactors_2_io_out_9_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_53_clock = clock;
  assign DFT_r_v2_53_reset = reset;
  assign DFT_r_v2_53_io_in_0_Re = TwiddleFactors_2_io_out_10_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_53_io_in_0_Im = TwiddleFactors_2_io_out_10_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_53_io_in_1_Re = TwiddleFactors_2_io_out_11_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_53_io_in_1_Im = TwiddleFactors_2_io_out_11_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_54_clock = clock;
  assign DFT_r_v2_54_reset = reset;
  assign DFT_r_v2_54_io_in_0_Re = TwiddleFactors_2_io_out_12_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_54_io_in_0_Im = TwiddleFactors_2_io_out_12_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_54_io_in_1_Re = TwiddleFactors_2_io_out_13_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_54_io_in_1_Im = TwiddleFactors_2_io_out_13_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_55_clock = clock;
  assign DFT_r_v2_55_reset = reset;
  assign DFT_r_v2_55_io_in_0_Re = TwiddleFactors_2_io_out_14_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_55_io_in_0_Im = TwiddleFactors_2_io_out_14_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_55_io_in_1_Re = TwiddleFactors_2_io_out_15_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_55_io_in_1_Im = TwiddleFactors_2_io_out_15_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_56_clock = clock;
  assign DFT_r_v2_56_reset = reset;
  assign DFT_r_v2_56_io_in_0_Re = TwiddleFactors_2_io_out_16_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_56_io_in_0_Im = TwiddleFactors_2_io_out_16_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_56_io_in_1_Re = TwiddleFactors_2_io_out_17_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_56_io_in_1_Im = TwiddleFactors_2_io_out_17_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_57_clock = clock;
  assign DFT_r_v2_57_reset = reset;
  assign DFT_r_v2_57_io_in_0_Re = TwiddleFactors_2_io_out_18_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_57_io_in_0_Im = TwiddleFactors_2_io_out_18_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_57_io_in_1_Re = TwiddleFactors_2_io_out_19_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_57_io_in_1_Im = TwiddleFactors_2_io_out_19_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_58_clock = clock;
  assign DFT_r_v2_58_reset = reset;
  assign DFT_r_v2_58_io_in_0_Re = TwiddleFactors_2_io_out_20_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_58_io_in_0_Im = TwiddleFactors_2_io_out_20_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_58_io_in_1_Re = TwiddleFactors_2_io_out_21_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_58_io_in_1_Im = TwiddleFactors_2_io_out_21_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_59_clock = clock;
  assign DFT_r_v2_59_reset = reset;
  assign DFT_r_v2_59_io_in_0_Re = TwiddleFactors_2_io_out_22_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_59_io_in_0_Im = TwiddleFactors_2_io_out_22_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_59_io_in_1_Re = TwiddleFactors_2_io_out_23_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_59_io_in_1_Im = TwiddleFactors_2_io_out_23_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_60_clock = clock;
  assign DFT_r_v2_60_reset = reset;
  assign DFT_r_v2_60_io_in_0_Re = TwiddleFactors_2_io_out_24_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_60_io_in_0_Im = TwiddleFactors_2_io_out_24_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_60_io_in_1_Re = TwiddleFactors_2_io_out_25_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_60_io_in_1_Im = TwiddleFactors_2_io_out_25_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_61_clock = clock;
  assign DFT_r_v2_61_reset = reset;
  assign DFT_r_v2_61_io_in_0_Re = TwiddleFactors_2_io_out_26_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_61_io_in_0_Im = TwiddleFactors_2_io_out_26_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_61_io_in_1_Re = TwiddleFactors_2_io_out_27_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_61_io_in_1_Im = TwiddleFactors_2_io_out_27_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_62_clock = clock;
  assign DFT_r_v2_62_reset = reset;
  assign DFT_r_v2_62_io_in_0_Re = TwiddleFactors_2_io_out_28_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_62_io_in_0_Im = TwiddleFactors_2_io_out_28_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_62_io_in_1_Re = TwiddleFactors_2_io_out_29_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_62_io_in_1_Im = TwiddleFactors_2_io_out_29_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_63_clock = clock;
  assign DFT_r_v2_63_reset = reset;
  assign DFT_r_v2_63_io_in_0_Re = TwiddleFactors_2_io_out_30_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_63_io_in_0_Im = TwiddleFactors_2_io_out_30_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_63_io_in_1_Re = TwiddleFactors_2_io_out_31_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_63_io_in_1_Im = TwiddleFactors_2_io_out_31_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_64_clock = clock;
  assign DFT_r_v2_64_reset = reset;
  assign DFT_r_v2_64_io_in_0_Re = TwiddleFactors_3_io_out_0_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_64_io_in_0_Im = TwiddleFactors_3_io_out_0_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_64_io_in_1_Re = TwiddleFactors_3_io_out_1_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_64_io_in_1_Im = TwiddleFactors_3_io_out_1_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_65_clock = clock;
  assign DFT_r_v2_65_reset = reset;
  assign DFT_r_v2_65_io_in_0_Re = TwiddleFactors_3_io_out_2_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_65_io_in_0_Im = TwiddleFactors_3_io_out_2_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_65_io_in_1_Re = TwiddleFactors_3_io_out_3_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_65_io_in_1_Im = TwiddleFactors_3_io_out_3_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_66_clock = clock;
  assign DFT_r_v2_66_reset = reset;
  assign DFT_r_v2_66_io_in_0_Re = TwiddleFactors_3_io_out_4_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_66_io_in_0_Im = TwiddleFactors_3_io_out_4_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_66_io_in_1_Re = TwiddleFactors_3_io_out_5_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_66_io_in_1_Im = TwiddleFactors_3_io_out_5_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_67_clock = clock;
  assign DFT_r_v2_67_reset = reset;
  assign DFT_r_v2_67_io_in_0_Re = TwiddleFactors_3_io_out_6_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_67_io_in_0_Im = TwiddleFactors_3_io_out_6_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_67_io_in_1_Re = TwiddleFactors_3_io_out_7_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_67_io_in_1_Im = TwiddleFactors_3_io_out_7_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_68_clock = clock;
  assign DFT_r_v2_68_reset = reset;
  assign DFT_r_v2_68_io_in_0_Re = TwiddleFactors_3_io_out_8_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_68_io_in_0_Im = TwiddleFactors_3_io_out_8_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_68_io_in_1_Re = TwiddleFactors_3_io_out_9_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_68_io_in_1_Im = TwiddleFactors_3_io_out_9_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_69_clock = clock;
  assign DFT_r_v2_69_reset = reset;
  assign DFT_r_v2_69_io_in_0_Re = TwiddleFactors_3_io_out_10_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_69_io_in_0_Im = TwiddleFactors_3_io_out_10_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_69_io_in_1_Re = TwiddleFactors_3_io_out_11_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_69_io_in_1_Im = TwiddleFactors_3_io_out_11_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_70_clock = clock;
  assign DFT_r_v2_70_reset = reset;
  assign DFT_r_v2_70_io_in_0_Re = TwiddleFactors_3_io_out_12_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_70_io_in_0_Im = TwiddleFactors_3_io_out_12_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_70_io_in_1_Re = TwiddleFactors_3_io_out_13_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_70_io_in_1_Im = TwiddleFactors_3_io_out_13_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_71_clock = clock;
  assign DFT_r_v2_71_reset = reset;
  assign DFT_r_v2_71_io_in_0_Re = TwiddleFactors_3_io_out_14_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_71_io_in_0_Im = TwiddleFactors_3_io_out_14_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_71_io_in_1_Re = TwiddleFactors_3_io_out_15_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_71_io_in_1_Im = TwiddleFactors_3_io_out_15_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_72_clock = clock;
  assign DFT_r_v2_72_reset = reset;
  assign DFT_r_v2_72_io_in_0_Re = TwiddleFactors_3_io_out_16_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_72_io_in_0_Im = TwiddleFactors_3_io_out_16_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_72_io_in_1_Re = TwiddleFactors_3_io_out_17_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_72_io_in_1_Im = TwiddleFactors_3_io_out_17_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_73_clock = clock;
  assign DFT_r_v2_73_reset = reset;
  assign DFT_r_v2_73_io_in_0_Re = TwiddleFactors_3_io_out_18_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_73_io_in_0_Im = TwiddleFactors_3_io_out_18_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_73_io_in_1_Re = TwiddleFactors_3_io_out_19_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_73_io_in_1_Im = TwiddleFactors_3_io_out_19_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_74_clock = clock;
  assign DFT_r_v2_74_reset = reset;
  assign DFT_r_v2_74_io_in_0_Re = TwiddleFactors_3_io_out_20_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_74_io_in_0_Im = TwiddleFactors_3_io_out_20_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_74_io_in_1_Re = TwiddleFactors_3_io_out_21_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_74_io_in_1_Im = TwiddleFactors_3_io_out_21_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_75_clock = clock;
  assign DFT_r_v2_75_reset = reset;
  assign DFT_r_v2_75_io_in_0_Re = TwiddleFactors_3_io_out_22_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_75_io_in_0_Im = TwiddleFactors_3_io_out_22_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_75_io_in_1_Re = TwiddleFactors_3_io_out_23_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_75_io_in_1_Im = TwiddleFactors_3_io_out_23_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_76_clock = clock;
  assign DFT_r_v2_76_reset = reset;
  assign DFT_r_v2_76_io_in_0_Re = TwiddleFactors_3_io_out_24_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_76_io_in_0_Im = TwiddleFactors_3_io_out_24_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_76_io_in_1_Re = TwiddleFactors_3_io_out_25_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_76_io_in_1_Im = TwiddleFactors_3_io_out_25_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_77_clock = clock;
  assign DFT_r_v2_77_reset = reset;
  assign DFT_r_v2_77_io_in_0_Re = TwiddleFactors_3_io_out_26_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_77_io_in_0_Im = TwiddleFactors_3_io_out_26_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_77_io_in_1_Re = TwiddleFactors_3_io_out_27_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_77_io_in_1_Im = TwiddleFactors_3_io_out_27_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_78_clock = clock;
  assign DFT_r_v2_78_reset = reset;
  assign DFT_r_v2_78_io_in_0_Re = TwiddleFactors_3_io_out_28_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_78_io_in_0_Im = TwiddleFactors_3_io_out_28_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_78_io_in_1_Re = TwiddleFactors_3_io_out_29_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_78_io_in_1_Im = TwiddleFactors_3_io_out_29_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_79_clock = clock;
  assign DFT_r_v2_79_reset = reset;
  assign DFT_r_v2_79_io_in_0_Re = TwiddleFactors_3_io_out_30_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_79_io_in_0_Im = TwiddleFactors_3_io_out_30_Im; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_79_io_in_1_Re = TwiddleFactors_3_io_out_31_Re; // @[FFTDesigns.scala 3147:39]
  assign DFT_r_v2_79_io_in_1_Im = TwiddleFactors_3_io_out_31_Im; // @[FFTDesigns.scala 3147:39]
  assign PermutationsBasic_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_2_Re = io_in_2_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_2_Im = io_in_2_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_3_Re = io_in_3_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_3_Im = io_in_3_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_4_Re = io_in_4_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_4_Im = io_in_4_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_5_Re = io_in_5_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_5_Im = io_in_5_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_6_Re = io_in_6_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_6_Im = io_in_6_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_7_Re = io_in_7_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_7_Im = io_in_7_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_8_Re = io_in_8_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_8_Im = io_in_8_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_9_Re = io_in_9_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_9_Im = io_in_9_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_10_Re = io_in_10_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_10_Im = io_in_10_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_11_Re = io_in_11_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_11_Im = io_in_11_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_12_Re = io_in_12_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_12_Im = io_in_12_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_13_Re = io_in_13_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_13_Im = io_in_13_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_14_Re = io_in_14_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_14_Im = io_in_14_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_15_Re = io_in_15_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_15_Im = io_in_15_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_16_Re = io_in_16_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_16_Im = io_in_16_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_17_Re = io_in_17_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_17_Im = io_in_17_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_18_Re = io_in_18_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_18_Im = io_in_18_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_19_Re = io_in_19_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_19_Im = io_in_19_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_20_Re = io_in_20_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_20_Im = io_in_20_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_21_Re = io_in_21_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_21_Im = io_in_21_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_22_Re = io_in_22_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_22_Im = io_in_22_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_23_Re = io_in_23_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_23_Im = io_in_23_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_24_Re = io_in_24_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_24_Im = io_in_24_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_25_Re = io_in_25_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_25_Im = io_in_25_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_26_Re = io_in_26_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_26_Im = io_in_26_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_27_Re = io_in_27_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_27_Im = io_in_27_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_28_Re = io_in_28_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_28_Im = io_in_28_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_29_Re = io_in_29_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_29_Im = io_in_29_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_30_Re = io_in_30_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_30_Im = io_in_30_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_31_Re = io_in_31_Re; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_io_in_31_Im = io_in_31_Im; // @[FFTDesigns.scala 3137:31]
  assign PermutationsBasic_1_io_in_0_Re = DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_0_Im = DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_1_Re = DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_1_Im = DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_2_Re = DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_2_Im = DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_3_Re = DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_3_Im = DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_4_Re = DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_4_Im = DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_5_Re = DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_5_Im = DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_6_Re = DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_6_Im = DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_7_Re = DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_7_Im = DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_8_Re = DFT_r_v2_4_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_8_Im = DFT_r_v2_4_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_9_Re = DFT_r_v2_4_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_9_Im = DFT_r_v2_4_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_10_Re = DFT_r_v2_5_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_10_Im = DFT_r_v2_5_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_11_Re = DFT_r_v2_5_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_11_Im = DFT_r_v2_5_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_12_Re = DFT_r_v2_6_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_12_Im = DFT_r_v2_6_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_13_Re = DFT_r_v2_6_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_13_Im = DFT_r_v2_6_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_14_Re = DFT_r_v2_7_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_14_Im = DFT_r_v2_7_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_15_Re = DFT_r_v2_7_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_15_Im = DFT_r_v2_7_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_16_Re = DFT_r_v2_8_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_16_Im = DFT_r_v2_8_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_17_Re = DFT_r_v2_8_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_17_Im = DFT_r_v2_8_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_18_Re = DFT_r_v2_9_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_18_Im = DFT_r_v2_9_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_19_Re = DFT_r_v2_9_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_19_Im = DFT_r_v2_9_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_20_Re = DFT_r_v2_10_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_20_Im = DFT_r_v2_10_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_21_Re = DFT_r_v2_10_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_21_Im = DFT_r_v2_10_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_22_Re = DFT_r_v2_11_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_22_Im = DFT_r_v2_11_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_23_Re = DFT_r_v2_11_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_23_Im = DFT_r_v2_11_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_24_Re = DFT_r_v2_12_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_24_Im = DFT_r_v2_12_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_25_Re = DFT_r_v2_12_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_25_Im = DFT_r_v2_12_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_26_Re = DFT_r_v2_13_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_26_Im = DFT_r_v2_13_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_27_Re = DFT_r_v2_13_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_27_Im = DFT_r_v2_13_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_28_Re = DFT_r_v2_14_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_28_Im = DFT_r_v2_14_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_29_Re = DFT_r_v2_14_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_29_Im = DFT_r_v2_14_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_30_Re = DFT_r_v2_15_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_30_Im = DFT_r_v2_15_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_31_Re = DFT_r_v2_15_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_1_io_in_31_Im = DFT_r_v2_15_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_0_Re = DFT_r_v2_16_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_0_Im = DFT_r_v2_16_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_1_Re = DFT_r_v2_16_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_1_Im = DFT_r_v2_16_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_2_Re = DFT_r_v2_17_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_2_Im = DFT_r_v2_17_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_3_Re = DFT_r_v2_17_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_3_Im = DFT_r_v2_17_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_4_Re = DFT_r_v2_18_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_4_Im = DFT_r_v2_18_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_5_Re = DFT_r_v2_18_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_5_Im = DFT_r_v2_18_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_6_Re = DFT_r_v2_19_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_6_Im = DFT_r_v2_19_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_7_Re = DFT_r_v2_19_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_7_Im = DFT_r_v2_19_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_8_Re = DFT_r_v2_20_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_8_Im = DFT_r_v2_20_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_9_Re = DFT_r_v2_20_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_9_Im = DFT_r_v2_20_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_10_Re = DFT_r_v2_21_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_10_Im = DFT_r_v2_21_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_11_Re = DFT_r_v2_21_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_11_Im = DFT_r_v2_21_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_12_Re = DFT_r_v2_22_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_12_Im = DFT_r_v2_22_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_13_Re = DFT_r_v2_22_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_13_Im = DFT_r_v2_22_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_14_Re = DFT_r_v2_23_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_14_Im = DFT_r_v2_23_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_15_Re = DFT_r_v2_23_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_15_Im = DFT_r_v2_23_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_16_Re = DFT_r_v2_24_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_16_Im = DFT_r_v2_24_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_17_Re = DFT_r_v2_24_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_17_Im = DFT_r_v2_24_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_18_Re = DFT_r_v2_25_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_18_Im = DFT_r_v2_25_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_19_Re = DFT_r_v2_25_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_19_Im = DFT_r_v2_25_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_20_Re = DFT_r_v2_26_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_20_Im = DFT_r_v2_26_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_21_Re = DFT_r_v2_26_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_21_Im = DFT_r_v2_26_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_22_Re = DFT_r_v2_27_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_22_Im = DFT_r_v2_27_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_23_Re = DFT_r_v2_27_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_23_Im = DFT_r_v2_27_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_24_Re = DFT_r_v2_28_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_24_Im = DFT_r_v2_28_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_25_Re = DFT_r_v2_28_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_25_Im = DFT_r_v2_28_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_26_Re = DFT_r_v2_29_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_26_Im = DFT_r_v2_29_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_27_Re = DFT_r_v2_29_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_27_Im = DFT_r_v2_29_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_28_Re = DFT_r_v2_30_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_28_Im = DFT_r_v2_30_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_29_Re = DFT_r_v2_30_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_29_Im = DFT_r_v2_30_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_30_Re = DFT_r_v2_31_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_30_Im = DFT_r_v2_31_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_31_Re = DFT_r_v2_31_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_2_io_in_31_Im = DFT_r_v2_31_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_0_Re = DFT_r_v2_32_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_0_Im = DFT_r_v2_32_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_1_Re = DFT_r_v2_32_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_1_Im = DFT_r_v2_32_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_2_Re = DFT_r_v2_33_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_2_Im = DFT_r_v2_33_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_3_Re = DFT_r_v2_33_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_3_Im = DFT_r_v2_33_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_4_Re = DFT_r_v2_34_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_4_Im = DFT_r_v2_34_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_5_Re = DFT_r_v2_34_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_5_Im = DFT_r_v2_34_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_6_Re = DFT_r_v2_35_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_6_Im = DFT_r_v2_35_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_7_Re = DFT_r_v2_35_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_7_Im = DFT_r_v2_35_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_8_Re = DFT_r_v2_36_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_8_Im = DFT_r_v2_36_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_9_Re = DFT_r_v2_36_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_9_Im = DFT_r_v2_36_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_10_Re = DFT_r_v2_37_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_10_Im = DFT_r_v2_37_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_11_Re = DFT_r_v2_37_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_11_Im = DFT_r_v2_37_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_12_Re = DFT_r_v2_38_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_12_Im = DFT_r_v2_38_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_13_Re = DFT_r_v2_38_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_13_Im = DFT_r_v2_38_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_14_Re = DFT_r_v2_39_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_14_Im = DFT_r_v2_39_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_15_Re = DFT_r_v2_39_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_15_Im = DFT_r_v2_39_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_16_Re = DFT_r_v2_40_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_16_Im = DFT_r_v2_40_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_17_Re = DFT_r_v2_40_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_17_Im = DFT_r_v2_40_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_18_Re = DFT_r_v2_41_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_18_Im = DFT_r_v2_41_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_19_Re = DFT_r_v2_41_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_19_Im = DFT_r_v2_41_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_20_Re = DFT_r_v2_42_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_20_Im = DFT_r_v2_42_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_21_Re = DFT_r_v2_42_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_21_Im = DFT_r_v2_42_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_22_Re = DFT_r_v2_43_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_22_Im = DFT_r_v2_43_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_23_Re = DFT_r_v2_43_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_23_Im = DFT_r_v2_43_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_24_Re = DFT_r_v2_44_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_24_Im = DFT_r_v2_44_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_25_Re = DFT_r_v2_44_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_25_Im = DFT_r_v2_44_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_26_Re = DFT_r_v2_45_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_26_Im = DFT_r_v2_45_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_27_Re = DFT_r_v2_45_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_27_Im = DFT_r_v2_45_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_28_Re = DFT_r_v2_46_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_28_Im = DFT_r_v2_46_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_29_Re = DFT_r_v2_46_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_29_Im = DFT_r_v2_46_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_30_Re = DFT_r_v2_47_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_30_Im = DFT_r_v2_47_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_31_Re = DFT_r_v2_47_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_3_io_in_31_Im = DFT_r_v2_47_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_0_Re = DFT_r_v2_48_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_0_Im = DFT_r_v2_48_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_1_Re = DFT_r_v2_48_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_1_Im = DFT_r_v2_48_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_2_Re = DFT_r_v2_49_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_2_Im = DFT_r_v2_49_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_3_Re = DFT_r_v2_49_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_3_Im = DFT_r_v2_49_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_4_Re = DFT_r_v2_50_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_4_Im = DFT_r_v2_50_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_5_Re = DFT_r_v2_50_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_5_Im = DFT_r_v2_50_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_6_Re = DFT_r_v2_51_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_6_Im = DFT_r_v2_51_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_7_Re = DFT_r_v2_51_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_7_Im = DFT_r_v2_51_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_8_Re = DFT_r_v2_52_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_8_Im = DFT_r_v2_52_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_9_Re = DFT_r_v2_52_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_9_Im = DFT_r_v2_52_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_10_Re = DFT_r_v2_53_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_10_Im = DFT_r_v2_53_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_11_Re = DFT_r_v2_53_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_11_Im = DFT_r_v2_53_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_12_Re = DFT_r_v2_54_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_12_Im = DFT_r_v2_54_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_13_Re = DFT_r_v2_54_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_13_Im = DFT_r_v2_54_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_14_Re = DFT_r_v2_55_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_14_Im = DFT_r_v2_55_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_15_Re = DFT_r_v2_55_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_15_Im = DFT_r_v2_55_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_16_Re = DFT_r_v2_56_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_16_Im = DFT_r_v2_56_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_17_Re = DFT_r_v2_56_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_17_Im = DFT_r_v2_56_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_18_Re = DFT_r_v2_57_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_18_Im = DFT_r_v2_57_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_19_Re = DFT_r_v2_57_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_19_Im = DFT_r_v2_57_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_20_Re = DFT_r_v2_58_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_20_Im = DFT_r_v2_58_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_21_Re = DFT_r_v2_58_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_21_Im = DFT_r_v2_58_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_22_Re = DFT_r_v2_59_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_22_Im = DFT_r_v2_59_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_23_Re = DFT_r_v2_59_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_23_Im = DFT_r_v2_59_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_24_Re = DFT_r_v2_60_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_24_Im = DFT_r_v2_60_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_25_Re = DFT_r_v2_60_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_25_Im = DFT_r_v2_60_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_26_Re = DFT_r_v2_61_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_26_Im = DFT_r_v2_61_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_27_Re = DFT_r_v2_61_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_27_Im = DFT_r_v2_61_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_28_Re = DFT_r_v2_62_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_28_Im = DFT_r_v2_62_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_29_Re = DFT_r_v2_62_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_29_Im = DFT_r_v2_62_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_30_Re = DFT_r_v2_63_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_30_Im = DFT_r_v2_63_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_31_Re = DFT_r_v2_63_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_4_io_in_31_Im = DFT_r_v2_63_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_0_Re = DFT_r_v2_64_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_0_Im = DFT_r_v2_64_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_1_Re = DFT_r_v2_64_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_1_Im = DFT_r_v2_64_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_2_Re = DFT_r_v2_65_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_2_Im = DFT_r_v2_65_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_3_Re = DFT_r_v2_65_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_3_Im = DFT_r_v2_65_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_4_Re = DFT_r_v2_66_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_4_Im = DFT_r_v2_66_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_5_Re = DFT_r_v2_66_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_5_Im = DFT_r_v2_66_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_6_Re = DFT_r_v2_67_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_6_Im = DFT_r_v2_67_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_7_Re = DFT_r_v2_67_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_7_Im = DFT_r_v2_67_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_8_Re = DFT_r_v2_68_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_8_Im = DFT_r_v2_68_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_9_Re = DFT_r_v2_68_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_9_Im = DFT_r_v2_68_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_10_Re = DFT_r_v2_69_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_10_Im = DFT_r_v2_69_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_11_Re = DFT_r_v2_69_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_11_Im = DFT_r_v2_69_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_12_Re = DFT_r_v2_70_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_12_Im = DFT_r_v2_70_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_13_Re = DFT_r_v2_70_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_13_Im = DFT_r_v2_70_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_14_Re = DFT_r_v2_71_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_14_Im = DFT_r_v2_71_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_15_Re = DFT_r_v2_71_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_15_Im = DFT_r_v2_71_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_16_Re = DFT_r_v2_72_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_16_Im = DFT_r_v2_72_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_17_Re = DFT_r_v2_72_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_17_Im = DFT_r_v2_72_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_18_Re = DFT_r_v2_73_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_18_Im = DFT_r_v2_73_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_19_Re = DFT_r_v2_73_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_19_Im = DFT_r_v2_73_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_20_Re = DFT_r_v2_74_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_20_Im = DFT_r_v2_74_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_21_Re = DFT_r_v2_74_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_21_Im = DFT_r_v2_74_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_22_Re = DFT_r_v2_75_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_22_Im = DFT_r_v2_75_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_23_Re = DFT_r_v2_75_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_23_Im = DFT_r_v2_75_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_24_Re = DFT_r_v2_76_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_24_Im = DFT_r_v2_76_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_25_Re = DFT_r_v2_76_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_25_Im = DFT_r_v2_76_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_26_Re = DFT_r_v2_77_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_26_Im = DFT_r_v2_77_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_27_Re = DFT_r_v2_77_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_27_Im = DFT_r_v2_77_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_28_Re = DFT_r_v2_78_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_28_Im = DFT_r_v2_78_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_29_Re = DFT_r_v2_78_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_29_Im = DFT_r_v2_78_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_30_Re = DFT_r_v2_79_io_out_0_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_30_Im = DFT_r_v2_79_io_out_0_Im; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_31_Re = DFT_r_v2_79_io_out_1_Re; // @[FFTDesigns.scala 3149:43]
  assign PermutationsBasic_5_io_in_31_Im = DFT_r_v2_79_io_out_1_Im; // @[FFTDesigns.scala 3149:43]
  assign TwiddleFactors_io_in_0_Re = PermutationsBasic_1_io_out_0_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_0_Im = PermutationsBasic_1_io_out_0_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_1_Re = PermutationsBasic_1_io_out_1_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_1_Im = PermutationsBasic_1_io_out_1_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_2_Re = PermutationsBasic_1_io_out_2_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_2_Im = PermutationsBasic_1_io_out_2_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_3_Re = PermutationsBasic_1_io_out_3_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_3_Im = PermutationsBasic_1_io_out_3_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_4_Re = PermutationsBasic_1_io_out_4_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_4_Im = PermutationsBasic_1_io_out_4_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_5_Re = PermutationsBasic_1_io_out_5_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_5_Im = PermutationsBasic_1_io_out_5_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_6_Re = PermutationsBasic_1_io_out_6_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_6_Im = PermutationsBasic_1_io_out_6_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_7_Re = PermutationsBasic_1_io_out_7_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_7_Im = PermutationsBasic_1_io_out_7_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_8_Re = PermutationsBasic_1_io_out_8_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_8_Im = PermutationsBasic_1_io_out_8_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_9_Re = PermutationsBasic_1_io_out_9_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_9_Im = PermutationsBasic_1_io_out_9_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_10_Re = PermutationsBasic_1_io_out_10_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_10_Im = PermutationsBasic_1_io_out_10_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_11_Re = PermutationsBasic_1_io_out_11_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_11_Im = PermutationsBasic_1_io_out_11_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_12_Re = PermutationsBasic_1_io_out_12_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_12_Im = PermutationsBasic_1_io_out_12_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_13_Re = PermutationsBasic_1_io_out_13_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_13_Im = PermutationsBasic_1_io_out_13_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_14_Re = PermutationsBasic_1_io_out_14_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_14_Im = PermutationsBasic_1_io_out_14_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_15_Re = PermutationsBasic_1_io_out_15_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_15_Im = PermutationsBasic_1_io_out_15_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_16_Re = PermutationsBasic_1_io_out_16_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_16_Im = PermutationsBasic_1_io_out_16_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_17_Re = PermutationsBasic_1_io_out_17_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_17_Im = PermutationsBasic_1_io_out_17_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_18_Re = PermutationsBasic_1_io_out_18_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_18_Im = PermutationsBasic_1_io_out_18_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_19_Re = PermutationsBasic_1_io_out_19_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_19_Im = PermutationsBasic_1_io_out_19_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_20_Re = PermutationsBasic_1_io_out_20_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_20_Im = PermutationsBasic_1_io_out_20_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_21_Re = PermutationsBasic_1_io_out_21_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_21_Im = PermutationsBasic_1_io_out_21_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_22_Re = PermutationsBasic_1_io_out_22_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_22_Im = PermutationsBasic_1_io_out_22_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_23_Re = PermutationsBasic_1_io_out_23_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_23_Im = PermutationsBasic_1_io_out_23_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_24_Re = PermutationsBasic_1_io_out_24_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_24_Im = PermutationsBasic_1_io_out_24_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_25_Re = PermutationsBasic_1_io_out_25_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_25_Im = PermutationsBasic_1_io_out_25_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_26_Re = PermutationsBasic_1_io_out_26_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_26_Im = PermutationsBasic_1_io_out_26_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_27_Re = PermutationsBasic_1_io_out_27_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_27_Im = PermutationsBasic_1_io_out_27_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_28_Re = PermutationsBasic_1_io_out_28_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_28_Im = PermutationsBasic_1_io_out_28_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_29_Re = PermutationsBasic_1_io_out_29_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_29_Im = PermutationsBasic_1_io_out_29_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_30_Re = PermutationsBasic_1_io_out_30_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_30_Im = PermutationsBasic_1_io_out_30_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_31_Re = PermutationsBasic_1_io_out_31_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_io_in_31_Im = PermutationsBasic_1_io_out_31_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_clock = clock;
  assign TwiddleFactors_1_reset = reset;
  assign TwiddleFactors_1_io_in_0_Re = PermutationsBasic_2_io_out_0_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_0_Im = PermutationsBasic_2_io_out_0_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_1_Re = PermutationsBasic_2_io_out_1_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_1_Im = PermutationsBasic_2_io_out_1_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_2_Re = PermutationsBasic_2_io_out_2_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_2_Im = PermutationsBasic_2_io_out_2_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_3_Re = PermutationsBasic_2_io_out_3_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_3_Im = PermutationsBasic_2_io_out_3_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_4_Re = PermutationsBasic_2_io_out_4_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_4_Im = PermutationsBasic_2_io_out_4_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_5_Re = PermutationsBasic_2_io_out_5_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_5_Im = PermutationsBasic_2_io_out_5_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_6_Re = PermutationsBasic_2_io_out_6_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_6_Im = PermutationsBasic_2_io_out_6_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_7_Re = PermutationsBasic_2_io_out_7_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_7_Im = PermutationsBasic_2_io_out_7_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_8_Re = PermutationsBasic_2_io_out_8_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_8_Im = PermutationsBasic_2_io_out_8_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_9_Re = PermutationsBasic_2_io_out_9_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_9_Im = PermutationsBasic_2_io_out_9_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_10_Re = PermutationsBasic_2_io_out_10_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_10_Im = PermutationsBasic_2_io_out_10_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_11_Re = PermutationsBasic_2_io_out_11_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_11_Im = PermutationsBasic_2_io_out_11_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_12_Re = PermutationsBasic_2_io_out_12_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_12_Im = PermutationsBasic_2_io_out_12_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_13_Re = PermutationsBasic_2_io_out_13_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_13_Im = PermutationsBasic_2_io_out_13_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_14_Re = PermutationsBasic_2_io_out_14_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_14_Im = PermutationsBasic_2_io_out_14_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_15_Re = PermutationsBasic_2_io_out_15_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_15_Im = PermutationsBasic_2_io_out_15_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_16_Re = PermutationsBasic_2_io_out_16_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_16_Im = PermutationsBasic_2_io_out_16_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_17_Re = PermutationsBasic_2_io_out_17_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_17_Im = PermutationsBasic_2_io_out_17_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_18_Re = PermutationsBasic_2_io_out_18_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_18_Im = PermutationsBasic_2_io_out_18_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_19_Re = PermutationsBasic_2_io_out_19_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_19_Im = PermutationsBasic_2_io_out_19_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_20_Re = PermutationsBasic_2_io_out_20_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_20_Im = PermutationsBasic_2_io_out_20_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_21_Re = PermutationsBasic_2_io_out_21_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_21_Im = PermutationsBasic_2_io_out_21_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_22_Re = PermutationsBasic_2_io_out_22_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_22_Im = PermutationsBasic_2_io_out_22_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_23_Re = PermutationsBasic_2_io_out_23_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_23_Im = PermutationsBasic_2_io_out_23_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_24_Re = PermutationsBasic_2_io_out_24_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_24_Im = PermutationsBasic_2_io_out_24_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_25_Re = PermutationsBasic_2_io_out_25_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_25_Im = PermutationsBasic_2_io_out_25_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_26_Re = PermutationsBasic_2_io_out_26_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_26_Im = PermutationsBasic_2_io_out_26_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_27_Re = PermutationsBasic_2_io_out_27_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_27_Im = PermutationsBasic_2_io_out_27_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_28_Re = PermutationsBasic_2_io_out_28_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_28_Im = PermutationsBasic_2_io_out_28_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_29_Re = PermutationsBasic_2_io_out_29_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_29_Im = PermutationsBasic_2_io_out_29_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_30_Re = PermutationsBasic_2_io_out_30_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_30_Im = PermutationsBasic_2_io_out_30_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_31_Re = PermutationsBasic_2_io_out_31_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_1_io_in_31_Im = PermutationsBasic_2_io_out_31_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_clock = clock;
  assign TwiddleFactors_2_reset = reset;
  assign TwiddleFactors_2_io_in_0_Re = PermutationsBasic_3_io_out_0_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_0_Im = PermutationsBasic_3_io_out_0_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_1_Re = PermutationsBasic_3_io_out_1_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_1_Im = PermutationsBasic_3_io_out_1_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_2_Re = PermutationsBasic_3_io_out_2_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_2_Im = PermutationsBasic_3_io_out_2_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_3_Re = PermutationsBasic_3_io_out_3_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_3_Im = PermutationsBasic_3_io_out_3_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_4_Re = PermutationsBasic_3_io_out_4_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_4_Im = PermutationsBasic_3_io_out_4_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_5_Re = PermutationsBasic_3_io_out_5_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_5_Im = PermutationsBasic_3_io_out_5_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_6_Re = PermutationsBasic_3_io_out_6_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_6_Im = PermutationsBasic_3_io_out_6_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_7_Re = PermutationsBasic_3_io_out_7_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_7_Im = PermutationsBasic_3_io_out_7_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_8_Re = PermutationsBasic_3_io_out_8_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_8_Im = PermutationsBasic_3_io_out_8_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_9_Re = PermutationsBasic_3_io_out_9_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_9_Im = PermutationsBasic_3_io_out_9_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_10_Re = PermutationsBasic_3_io_out_10_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_10_Im = PermutationsBasic_3_io_out_10_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_11_Re = PermutationsBasic_3_io_out_11_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_11_Im = PermutationsBasic_3_io_out_11_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_12_Re = PermutationsBasic_3_io_out_12_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_12_Im = PermutationsBasic_3_io_out_12_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_13_Re = PermutationsBasic_3_io_out_13_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_13_Im = PermutationsBasic_3_io_out_13_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_14_Re = PermutationsBasic_3_io_out_14_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_14_Im = PermutationsBasic_3_io_out_14_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_15_Re = PermutationsBasic_3_io_out_15_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_15_Im = PermutationsBasic_3_io_out_15_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_16_Re = PermutationsBasic_3_io_out_16_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_16_Im = PermutationsBasic_3_io_out_16_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_17_Re = PermutationsBasic_3_io_out_17_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_17_Im = PermutationsBasic_3_io_out_17_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_18_Re = PermutationsBasic_3_io_out_18_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_18_Im = PermutationsBasic_3_io_out_18_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_19_Re = PermutationsBasic_3_io_out_19_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_19_Im = PermutationsBasic_3_io_out_19_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_20_Re = PermutationsBasic_3_io_out_20_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_20_Im = PermutationsBasic_3_io_out_20_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_21_Re = PermutationsBasic_3_io_out_21_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_21_Im = PermutationsBasic_3_io_out_21_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_22_Re = PermutationsBasic_3_io_out_22_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_22_Im = PermutationsBasic_3_io_out_22_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_23_Re = PermutationsBasic_3_io_out_23_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_23_Im = PermutationsBasic_3_io_out_23_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_24_Re = PermutationsBasic_3_io_out_24_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_24_Im = PermutationsBasic_3_io_out_24_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_25_Re = PermutationsBasic_3_io_out_25_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_25_Im = PermutationsBasic_3_io_out_25_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_26_Re = PermutationsBasic_3_io_out_26_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_26_Im = PermutationsBasic_3_io_out_26_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_27_Re = PermutationsBasic_3_io_out_27_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_27_Im = PermutationsBasic_3_io_out_27_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_28_Re = PermutationsBasic_3_io_out_28_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_28_Im = PermutationsBasic_3_io_out_28_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_29_Re = PermutationsBasic_3_io_out_29_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_29_Im = PermutationsBasic_3_io_out_29_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_30_Re = PermutationsBasic_3_io_out_30_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_30_Im = PermutationsBasic_3_io_out_30_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_31_Re = PermutationsBasic_3_io_out_31_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_2_io_in_31_Im = PermutationsBasic_3_io_out_31_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_clock = clock;
  assign TwiddleFactors_3_reset = reset;
  assign TwiddleFactors_3_io_in_0_Re = PermutationsBasic_4_io_out_0_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_0_Im = PermutationsBasic_4_io_out_0_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_1_Re = PermutationsBasic_4_io_out_1_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_1_Im = PermutationsBasic_4_io_out_1_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_2_Re = PermutationsBasic_4_io_out_2_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_2_Im = PermutationsBasic_4_io_out_2_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_3_Re = PermutationsBasic_4_io_out_3_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_3_Im = PermutationsBasic_4_io_out_3_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_4_Re = PermutationsBasic_4_io_out_4_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_4_Im = PermutationsBasic_4_io_out_4_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_5_Re = PermutationsBasic_4_io_out_5_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_5_Im = PermutationsBasic_4_io_out_5_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_6_Re = PermutationsBasic_4_io_out_6_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_6_Im = PermutationsBasic_4_io_out_6_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_7_Re = PermutationsBasic_4_io_out_7_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_7_Im = PermutationsBasic_4_io_out_7_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_8_Re = PermutationsBasic_4_io_out_8_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_8_Im = PermutationsBasic_4_io_out_8_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_9_Re = PermutationsBasic_4_io_out_9_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_9_Im = PermutationsBasic_4_io_out_9_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_10_Re = PermutationsBasic_4_io_out_10_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_10_Im = PermutationsBasic_4_io_out_10_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_11_Re = PermutationsBasic_4_io_out_11_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_11_Im = PermutationsBasic_4_io_out_11_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_12_Re = PermutationsBasic_4_io_out_12_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_12_Im = PermutationsBasic_4_io_out_12_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_13_Re = PermutationsBasic_4_io_out_13_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_13_Im = PermutationsBasic_4_io_out_13_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_14_Re = PermutationsBasic_4_io_out_14_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_14_Im = PermutationsBasic_4_io_out_14_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_15_Re = PermutationsBasic_4_io_out_15_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_15_Im = PermutationsBasic_4_io_out_15_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_16_Re = PermutationsBasic_4_io_out_16_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_16_Im = PermutationsBasic_4_io_out_16_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_17_Re = PermutationsBasic_4_io_out_17_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_17_Im = PermutationsBasic_4_io_out_17_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_18_Re = PermutationsBasic_4_io_out_18_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_18_Im = PermutationsBasic_4_io_out_18_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_19_Re = PermutationsBasic_4_io_out_19_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_19_Im = PermutationsBasic_4_io_out_19_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_20_Re = PermutationsBasic_4_io_out_20_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_20_Im = PermutationsBasic_4_io_out_20_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_21_Re = PermutationsBasic_4_io_out_21_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_21_Im = PermutationsBasic_4_io_out_21_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_22_Re = PermutationsBasic_4_io_out_22_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_22_Im = PermutationsBasic_4_io_out_22_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_23_Re = PermutationsBasic_4_io_out_23_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_23_Im = PermutationsBasic_4_io_out_23_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_24_Re = PermutationsBasic_4_io_out_24_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_24_Im = PermutationsBasic_4_io_out_24_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_25_Re = PermutationsBasic_4_io_out_25_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_25_Im = PermutationsBasic_4_io_out_25_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_26_Re = PermutationsBasic_4_io_out_26_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_26_Im = PermutationsBasic_4_io_out_26_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_27_Re = PermutationsBasic_4_io_out_27_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_27_Im = PermutationsBasic_4_io_out_27_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_28_Re = PermutationsBasic_4_io_out_28_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_28_Im = PermutationsBasic_4_io_out_28_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_29_Re = PermutationsBasic_4_io_out_29_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_29_Im = PermutationsBasic_4_io_out_29_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_30_Re = PermutationsBasic_4_io_out_30_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_30_Im = PermutationsBasic_4_io_out_30_Im; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_31_Re = PermutationsBasic_4_io_out_31_Re; // @[FFTDesigns.scala 3153:38]
  assign TwiddleFactors_3_io_in_31_Im = PermutationsBasic_4_io_out_31_Im; // @[FFTDesigns.scala 3153:38]
endmodule
module PermutationsBasic_82(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  input  [31:0] io_in_32_Re,
  input  [31:0] io_in_32_Im,
  input  [31:0] io_in_33_Re,
  input  [31:0] io_in_33_Im,
  input  [31:0] io_in_34_Re,
  input  [31:0] io_in_34_Im,
  input  [31:0] io_in_35_Re,
  input  [31:0] io_in_35_Im,
  input  [31:0] io_in_36_Re,
  input  [31:0] io_in_36_Im,
  input  [31:0] io_in_37_Re,
  input  [31:0] io_in_37_Im,
  input  [31:0] io_in_38_Re,
  input  [31:0] io_in_38_Im,
  input  [31:0] io_in_39_Re,
  input  [31:0] io_in_39_Im,
  input  [31:0] io_in_40_Re,
  input  [31:0] io_in_40_Im,
  input  [31:0] io_in_41_Re,
  input  [31:0] io_in_41_Im,
  input  [31:0] io_in_42_Re,
  input  [31:0] io_in_42_Im,
  input  [31:0] io_in_43_Re,
  input  [31:0] io_in_43_Im,
  input  [31:0] io_in_44_Re,
  input  [31:0] io_in_44_Im,
  input  [31:0] io_in_45_Re,
  input  [31:0] io_in_45_Im,
  input  [31:0] io_in_46_Re,
  input  [31:0] io_in_46_Im,
  input  [31:0] io_in_47_Re,
  input  [31:0] io_in_47_Im,
  input  [31:0] io_in_48_Re,
  input  [31:0] io_in_48_Im,
  input  [31:0] io_in_49_Re,
  input  [31:0] io_in_49_Im,
  input  [31:0] io_in_50_Re,
  input  [31:0] io_in_50_Im,
  input  [31:0] io_in_51_Re,
  input  [31:0] io_in_51_Im,
  input  [31:0] io_in_52_Re,
  input  [31:0] io_in_52_Im,
  input  [31:0] io_in_53_Re,
  input  [31:0] io_in_53_Im,
  input  [31:0] io_in_54_Re,
  input  [31:0] io_in_54_Im,
  input  [31:0] io_in_55_Re,
  input  [31:0] io_in_55_Im,
  input  [31:0] io_in_56_Re,
  input  [31:0] io_in_56_Im,
  input  [31:0] io_in_57_Re,
  input  [31:0] io_in_57_Im,
  input  [31:0] io_in_58_Re,
  input  [31:0] io_in_58_Im,
  input  [31:0] io_in_59_Re,
  input  [31:0] io_in_59_Im,
  input  [31:0] io_in_60_Re,
  input  [31:0] io_in_60_Im,
  input  [31:0] io_in_61_Re,
  input  [31:0] io_in_61_Im,
  input  [31:0] io_in_62_Re,
  input  [31:0] io_in_62_Im,
  input  [31:0] io_in_63_Re,
  input  [31:0] io_in_63_Im,
  input  [31:0] io_in_64_Re,
  input  [31:0] io_in_64_Im,
  input  [31:0] io_in_65_Re,
  input  [31:0] io_in_65_Im,
  input  [31:0] io_in_66_Re,
  input  [31:0] io_in_66_Im,
  input  [31:0] io_in_67_Re,
  input  [31:0] io_in_67_Im,
  input  [31:0] io_in_68_Re,
  input  [31:0] io_in_68_Im,
  input  [31:0] io_in_69_Re,
  input  [31:0] io_in_69_Im,
  input  [31:0] io_in_70_Re,
  input  [31:0] io_in_70_Im,
  input  [31:0] io_in_71_Re,
  input  [31:0] io_in_71_Im,
  input  [31:0] io_in_72_Re,
  input  [31:0] io_in_72_Im,
  input  [31:0] io_in_73_Re,
  input  [31:0] io_in_73_Im,
  input  [31:0] io_in_74_Re,
  input  [31:0] io_in_74_Im,
  input  [31:0] io_in_75_Re,
  input  [31:0] io_in_75_Im,
  input  [31:0] io_in_76_Re,
  input  [31:0] io_in_76_Im,
  input  [31:0] io_in_77_Re,
  input  [31:0] io_in_77_Im,
  input  [31:0] io_in_78_Re,
  input  [31:0] io_in_78_Im,
  input  [31:0] io_in_79_Re,
  input  [31:0] io_in_79_Im,
  input  [31:0] io_in_80_Re,
  input  [31:0] io_in_80_Im,
  input  [31:0] io_in_81_Re,
  input  [31:0] io_in_81_Im,
  input  [31:0] io_in_82_Re,
  input  [31:0] io_in_82_Im,
  input  [31:0] io_in_83_Re,
  input  [31:0] io_in_83_Im,
  input  [31:0] io_in_84_Re,
  input  [31:0] io_in_84_Im,
  input  [31:0] io_in_85_Re,
  input  [31:0] io_in_85_Im,
  input  [31:0] io_in_86_Re,
  input  [31:0] io_in_86_Im,
  input  [31:0] io_in_87_Re,
  input  [31:0] io_in_87_Im,
  input  [31:0] io_in_88_Re,
  input  [31:0] io_in_88_Im,
  input  [31:0] io_in_89_Re,
  input  [31:0] io_in_89_Im,
  input  [31:0] io_in_90_Re,
  input  [31:0] io_in_90_Im,
  input  [31:0] io_in_91_Re,
  input  [31:0] io_in_91_Im,
  input  [31:0] io_in_92_Re,
  input  [31:0] io_in_92_Im,
  input  [31:0] io_in_93_Re,
  input  [31:0] io_in_93_Im,
  input  [31:0] io_in_94_Re,
  input  [31:0] io_in_94_Im,
  input  [31:0] io_in_95_Re,
  input  [31:0] io_in_95_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im,
  output [31:0] io_out_32_Re,
  output [31:0] io_out_32_Im,
  output [31:0] io_out_33_Re,
  output [31:0] io_out_33_Im,
  output [31:0] io_out_34_Re,
  output [31:0] io_out_34_Im,
  output [31:0] io_out_35_Re,
  output [31:0] io_out_35_Im,
  output [31:0] io_out_36_Re,
  output [31:0] io_out_36_Im,
  output [31:0] io_out_37_Re,
  output [31:0] io_out_37_Im,
  output [31:0] io_out_38_Re,
  output [31:0] io_out_38_Im,
  output [31:0] io_out_39_Re,
  output [31:0] io_out_39_Im,
  output [31:0] io_out_40_Re,
  output [31:0] io_out_40_Im,
  output [31:0] io_out_41_Re,
  output [31:0] io_out_41_Im,
  output [31:0] io_out_42_Re,
  output [31:0] io_out_42_Im,
  output [31:0] io_out_43_Re,
  output [31:0] io_out_43_Im,
  output [31:0] io_out_44_Re,
  output [31:0] io_out_44_Im,
  output [31:0] io_out_45_Re,
  output [31:0] io_out_45_Im,
  output [31:0] io_out_46_Re,
  output [31:0] io_out_46_Im,
  output [31:0] io_out_47_Re,
  output [31:0] io_out_47_Im,
  output [31:0] io_out_48_Re,
  output [31:0] io_out_48_Im,
  output [31:0] io_out_49_Re,
  output [31:0] io_out_49_Im,
  output [31:0] io_out_50_Re,
  output [31:0] io_out_50_Im,
  output [31:0] io_out_51_Re,
  output [31:0] io_out_51_Im,
  output [31:0] io_out_52_Re,
  output [31:0] io_out_52_Im,
  output [31:0] io_out_53_Re,
  output [31:0] io_out_53_Im,
  output [31:0] io_out_54_Re,
  output [31:0] io_out_54_Im,
  output [31:0] io_out_55_Re,
  output [31:0] io_out_55_Im,
  output [31:0] io_out_56_Re,
  output [31:0] io_out_56_Im,
  output [31:0] io_out_57_Re,
  output [31:0] io_out_57_Im,
  output [31:0] io_out_58_Re,
  output [31:0] io_out_58_Im,
  output [31:0] io_out_59_Re,
  output [31:0] io_out_59_Im,
  output [31:0] io_out_60_Re,
  output [31:0] io_out_60_Im,
  output [31:0] io_out_61_Re,
  output [31:0] io_out_61_Im,
  output [31:0] io_out_62_Re,
  output [31:0] io_out_62_Im,
  output [31:0] io_out_63_Re,
  output [31:0] io_out_63_Im,
  output [31:0] io_out_64_Re,
  output [31:0] io_out_64_Im,
  output [31:0] io_out_65_Re,
  output [31:0] io_out_65_Im,
  output [31:0] io_out_66_Re,
  output [31:0] io_out_66_Im,
  output [31:0] io_out_67_Re,
  output [31:0] io_out_67_Im,
  output [31:0] io_out_68_Re,
  output [31:0] io_out_68_Im,
  output [31:0] io_out_69_Re,
  output [31:0] io_out_69_Im,
  output [31:0] io_out_70_Re,
  output [31:0] io_out_70_Im,
  output [31:0] io_out_71_Re,
  output [31:0] io_out_71_Im,
  output [31:0] io_out_72_Re,
  output [31:0] io_out_72_Im,
  output [31:0] io_out_73_Re,
  output [31:0] io_out_73_Im,
  output [31:0] io_out_74_Re,
  output [31:0] io_out_74_Im,
  output [31:0] io_out_75_Re,
  output [31:0] io_out_75_Im,
  output [31:0] io_out_76_Re,
  output [31:0] io_out_76_Im,
  output [31:0] io_out_77_Re,
  output [31:0] io_out_77_Im,
  output [31:0] io_out_78_Re,
  output [31:0] io_out_78_Im,
  output [31:0] io_out_79_Re,
  output [31:0] io_out_79_Im,
  output [31:0] io_out_80_Re,
  output [31:0] io_out_80_Im,
  output [31:0] io_out_81_Re,
  output [31:0] io_out_81_Im,
  output [31:0] io_out_82_Re,
  output [31:0] io_out_82_Im,
  output [31:0] io_out_83_Re,
  output [31:0] io_out_83_Im,
  output [31:0] io_out_84_Re,
  output [31:0] io_out_84_Im,
  output [31:0] io_out_85_Re,
  output [31:0] io_out_85_Im,
  output [31:0] io_out_86_Re,
  output [31:0] io_out_86_Im,
  output [31:0] io_out_87_Re,
  output [31:0] io_out_87_Im,
  output [31:0] io_out_88_Re,
  output [31:0] io_out_88_Im,
  output [31:0] io_out_89_Re,
  output [31:0] io_out_89_Im,
  output [31:0] io_out_90_Re,
  output [31:0] io_out_90_Im,
  output [31:0] io_out_91_Re,
  output [31:0] io_out_91_Im,
  output [31:0] io_out_92_Re,
  output [31:0] io_out_92_Im,
  output [31:0] io_out_93_Re,
  output [31:0] io_out_93_Im,
  output [31:0] io_out_94_Re,
  output [31:0] io_out_94_Im,
  output [31:0] io_out_95_Re,
  output [31:0] io_out_95_Im
);
  assign io_out_0_Re = io_in_0_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_0_Im = io_in_0_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Re = io_in_32_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Im = io_in_32_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Re = io_in_64_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Im = io_in_64_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_3_Re = io_in_1_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_3_Im = io_in_1_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_4_Re = io_in_33_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_4_Im = io_in_33_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_5_Re = io_in_65_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_5_Im = io_in_65_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_6_Re = io_in_2_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_6_Im = io_in_2_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_7_Re = io_in_34_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_7_Im = io_in_34_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_8_Re = io_in_66_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_8_Im = io_in_66_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_9_Re = io_in_3_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_9_Im = io_in_3_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_10_Re = io_in_35_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_10_Im = io_in_35_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_11_Re = io_in_67_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_11_Im = io_in_67_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_12_Re = io_in_4_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_12_Im = io_in_4_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_13_Re = io_in_36_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_13_Im = io_in_36_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_14_Re = io_in_68_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_14_Im = io_in_68_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_15_Re = io_in_5_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_15_Im = io_in_5_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_16_Re = io_in_37_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_16_Im = io_in_37_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_17_Re = io_in_69_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_17_Im = io_in_69_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_18_Re = io_in_6_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_18_Im = io_in_6_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_19_Re = io_in_38_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_19_Im = io_in_38_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_20_Re = io_in_70_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_20_Im = io_in_70_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_21_Re = io_in_7_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_21_Im = io_in_7_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_22_Re = io_in_39_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_22_Im = io_in_39_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_23_Re = io_in_71_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_23_Im = io_in_71_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_24_Re = io_in_8_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_24_Im = io_in_8_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_25_Re = io_in_40_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_25_Im = io_in_40_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_26_Re = io_in_72_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_26_Im = io_in_72_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_27_Re = io_in_9_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_27_Im = io_in_9_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_28_Re = io_in_41_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_28_Im = io_in_41_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_29_Re = io_in_73_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_29_Im = io_in_73_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_30_Re = io_in_10_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_30_Im = io_in_10_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_31_Re = io_in_42_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_31_Im = io_in_42_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_32_Re = io_in_74_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_32_Im = io_in_74_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_33_Re = io_in_11_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_33_Im = io_in_11_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_34_Re = io_in_43_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_34_Im = io_in_43_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_35_Re = io_in_75_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_35_Im = io_in_75_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_36_Re = io_in_12_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_36_Im = io_in_12_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_37_Re = io_in_44_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_37_Im = io_in_44_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_38_Re = io_in_76_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_38_Im = io_in_76_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_39_Re = io_in_13_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_39_Im = io_in_13_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_40_Re = io_in_45_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_40_Im = io_in_45_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_41_Re = io_in_77_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_41_Im = io_in_77_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_42_Re = io_in_14_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_42_Im = io_in_14_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_43_Re = io_in_46_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_43_Im = io_in_46_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_44_Re = io_in_78_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_44_Im = io_in_78_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_45_Re = io_in_15_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_45_Im = io_in_15_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_46_Re = io_in_47_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_46_Im = io_in_47_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_47_Re = io_in_79_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_47_Im = io_in_79_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_48_Re = io_in_16_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_48_Im = io_in_16_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_49_Re = io_in_48_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_49_Im = io_in_48_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_50_Re = io_in_80_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_50_Im = io_in_80_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_51_Re = io_in_17_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_51_Im = io_in_17_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_52_Re = io_in_49_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_52_Im = io_in_49_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_53_Re = io_in_81_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_53_Im = io_in_81_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_54_Re = io_in_18_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_54_Im = io_in_18_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_55_Re = io_in_50_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_55_Im = io_in_50_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_56_Re = io_in_82_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_56_Im = io_in_82_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_57_Re = io_in_19_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_57_Im = io_in_19_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_58_Re = io_in_51_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_58_Im = io_in_51_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_59_Re = io_in_83_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_59_Im = io_in_83_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_60_Re = io_in_20_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_60_Im = io_in_20_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_61_Re = io_in_52_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_61_Im = io_in_52_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_62_Re = io_in_84_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_62_Im = io_in_84_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_63_Re = io_in_21_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_63_Im = io_in_21_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_64_Re = io_in_53_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_64_Im = io_in_53_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_65_Re = io_in_85_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_65_Im = io_in_85_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_66_Re = io_in_22_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_66_Im = io_in_22_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_67_Re = io_in_54_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_67_Im = io_in_54_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_68_Re = io_in_86_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_68_Im = io_in_86_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_69_Re = io_in_23_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_69_Im = io_in_23_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_70_Re = io_in_55_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_70_Im = io_in_55_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_71_Re = io_in_87_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_71_Im = io_in_87_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_72_Re = io_in_24_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_72_Im = io_in_24_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_73_Re = io_in_56_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_73_Im = io_in_56_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_74_Re = io_in_88_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_74_Im = io_in_88_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_75_Re = io_in_25_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_75_Im = io_in_25_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_76_Re = io_in_57_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_76_Im = io_in_57_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_77_Re = io_in_89_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_77_Im = io_in_89_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_78_Re = io_in_26_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_78_Im = io_in_26_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_79_Re = io_in_58_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_79_Im = io_in_58_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_80_Re = io_in_90_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_80_Im = io_in_90_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_81_Re = io_in_27_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_81_Im = io_in_27_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_82_Re = io_in_59_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_82_Im = io_in_59_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_83_Re = io_in_91_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_83_Im = io_in_91_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_84_Re = io_in_28_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_84_Im = io_in_28_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_85_Re = io_in_60_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_85_Im = io_in_60_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_86_Re = io_in_92_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_86_Im = io_in_92_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_87_Re = io_in_29_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_87_Im = io_in_29_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_88_Re = io_in_61_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_88_Im = io_in_61_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_89_Re = io_in_93_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_89_Im = io_in_93_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_90_Re = io_in_30_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_90_Im = io_in_30_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_91_Re = io_in_62_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_91_Im = io_in_62_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_92_Re = io_in_94_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_92_Im = io_in_94_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_93_Re = io_in_31_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_93_Im = io_in_31_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_94_Re = io_in_63_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_94_Im = io_in_63_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_95_Re = io_in_95_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_95_Im = io_in_95_Im; // @[FFTDesigns.scala 2315:17]
endmodule
module PermutationsBasic_83(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  input  [31:0] io_in_32_Re,
  input  [31:0] io_in_32_Im,
  input  [31:0] io_in_33_Re,
  input  [31:0] io_in_33_Im,
  input  [31:0] io_in_34_Re,
  input  [31:0] io_in_34_Im,
  input  [31:0] io_in_35_Re,
  input  [31:0] io_in_35_Im,
  input  [31:0] io_in_36_Re,
  input  [31:0] io_in_36_Im,
  input  [31:0] io_in_37_Re,
  input  [31:0] io_in_37_Im,
  input  [31:0] io_in_38_Re,
  input  [31:0] io_in_38_Im,
  input  [31:0] io_in_39_Re,
  input  [31:0] io_in_39_Im,
  input  [31:0] io_in_40_Re,
  input  [31:0] io_in_40_Im,
  input  [31:0] io_in_41_Re,
  input  [31:0] io_in_41_Im,
  input  [31:0] io_in_42_Re,
  input  [31:0] io_in_42_Im,
  input  [31:0] io_in_43_Re,
  input  [31:0] io_in_43_Im,
  input  [31:0] io_in_44_Re,
  input  [31:0] io_in_44_Im,
  input  [31:0] io_in_45_Re,
  input  [31:0] io_in_45_Im,
  input  [31:0] io_in_46_Re,
  input  [31:0] io_in_46_Im,
  input  [31:0] io_in_47_Re,
  input  [31:0] io_in_47_Im,
  input  [31:0] io_in_48_Re,
  input  [31:0] io_in_48_Im,
  input  [31:0] io_in_49_Re,
  input  [31:0] io_in_49_Im,
  input  [31:0] io_in_50_Re,
  input  [31:0] io_in_50_Im,
  input  [31:0] io_in_51_Re,
  input  [31:0] io_in_51_Im,
  input  [31:0] io_in_52_Re,
  input  [31:0] io_in_52_Im,
  input  [31:0] io_in_53_Re,
  input  [31:0] io_in_53_Im,
  input  [31:0] io_in_54_Re,
  input  [31:0] io_in_54_Im,
  input  [31:0] io_in_55_Re,
  input  [31:0] io_in_55_Im,
  input  [31:0] io_in_56_Re,
  input  [31:0] io_in_56_Im,
  input  [31:0] io_in_57_Re,
  input  [31:0] io_in_57_Im,
  input  [31:0] io_in_58_Re,
  input  [31:0] io_in_58_Im,
  input  [31:0] io_in_59_Re,
  input  [31:0] io_in_59_Im,
  input  [31:0] io_in_60_Re,
  input  [31:0] io_in_60_Im,
  input  [31:0] io_in_61_Re,
  input  [31:0] io_in_61_Im,
  input  [31:0] io_in_62_Re,
  input  [31:0] io_in_62_Im,
  input  [31:0] io_in_63_Re,
  input  [31:0] io_in_63_Im,
  input  [31:0] io_in_64_Re,
  input  [31:0] io_in_64_Im,
  input  [31:0] io_in_65_Re,
  input  [31:0] io_in_65_Im,
  input  [31:0] io_in_66_Re,
  input  [31:0] io_in_66_Im,
  input  [31:0] io_in_67_Re,
  input  [31:0] io_in_67_Im,
  input  [31:0] io_in_68_Re,
  input  [31:0] io_in_68_Im,
  input  [31:0] io_in_69_Re,
  input  [31:0] io_in_69_Im,
  input  [31:0] io_in_70_Re,
  input  [31:0] io_in_70_Im,
  input  [31:0] io_in_71_Re,
  input  [31:0] io_in_71_Im,
  input  [31:0] io_in_72_Re,
  input  [31:0] io_in_72_Im,
  input  [31:0] io_in_73_Re,
  input  [31:0] io_in_73_Im,
  input  [31:0] io_in_74_Re,
  input  [31:0] io_in_74_Im,
  input  [31:0] io_in_75_Re,
  input  [31:0] io_in_75_Im,
  input  [31:0] io_in_76_Re,
  input  [31:0] io_in_76_Im,
  input  [31:0] io_in_77_Re,
  input  [31:0] io_in_77_Im,
  input  [31:0] io_in_78_Re,
  input  [31:0] io_in_78_Im,
  input  [31:0] io_in_79_Re,
  input  [31:0] io_in_79_Im,
  input  [31:0] io_in_80_Re,
  input  [31:0] io_in_80_Im,
  input  [31:0] io_in_81_Re,
  input  [31:0] io_in_81_Im,
  input  [31:0] io_in_82_Re,
  input  [31:0] io_in_82_Im,
  input  [31:0] io_in_83_Re,
  input  [31:0] io_in_83_Im,
  input  [31:0] io_in_84_Re,
  input  [31:0] io_in_84_Im,
  input  [31:0] io_in_85_Re,
  input  [31:0] io_in_85_Im,
  input  [31:0] io_in_86_Re,
  input  [31:0] io_in_86_Im,
  input  [31:0] io_in_87_Re,
  input  [31:0] io_in_87_Im,
  input  [31:0] io_in_88_Re,
  input  [31:0] io_in_88_Im,
  input  [31:0] io_in_89_Re,
  input  [31:0] io_in_89_Im,
  input  [31:0] io_in_90_Re,
  input  [31:0] io_in_90_Im,
  input  [31:0] io_in_91_Re,
  input  [31:0] io_in_91_Im,
  input  [31:0] io_in_92_Re,
  input  [31:0] io_in_92_Im,
  input  [31:0] io_in_93_Re,
  input  [31:0] io_in_93_Im,
  input  [31:0] io_in_94_Re,
  input  [31:0] io_in_94_Im,
  input  [31:0] io_in_95_Re,
  input  [31:0] io_in_95_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im,
  output [31:0] io_out_32_Re,
  output [31:0] io_out_32_Im,
  output [31:0] io_out_33_Re,
  output [31:0] io_out_33_Im,
  output [31:0] io_out_34_Re,
  output [31:0] io_out_34_Im,
  output [31:0] io_out_35_Re,
  output [31:0] io_out_35_Im,
  output [31:0] io_out_36_Re,
  output [31:0] io_out_36_Im,
  output [31:0] io_out_37_Re,
  output [31:0] io_out_37_Im,
  output [31:0] io_out_38_Re,
  output [31:0] io_out_38_Im,
  output [31:0] io_out_39_Re,
  output [31:0] io_out_39_Im,
  output [31:0] io_out_40_Re,
  output [31:0] io_out_40_Im,
  output [31:0] io_out_41_Re,
  output [31:0] io_out_41_Im,
  output [31:0] io_out_42_Re,
  output [31:0] io_out_42_Im,
  output [31:0] io_out_43_Re,
  output [31:0] io_out_43_Im,
  output [31:0] io_out_44_Re,
  output [31:0] io_out_44_Im,
  output [31:0] io_out_45_Re,
  output [31:0] io_out_45_Im,
  output [31:0] io_out_46_Re,
  output [31:0] io_out_46_Im,
  output [31:0] io_out_47_Re,
  output [31:0] io_out_47_Im,
  output [31:0] io_out_48_Re,
  output [31:0] io_out_48_Im,
  output [31:0] io_out_49_Re,
  output [31:0] io_out_49_Im,
  output [31:0] io_out_50_Re,
  output [31:0] io_out_50_Im,
  output [31:0] io_out_51_Re,
  output [31:0] io_out_51_Im,
  output [31:0] io_out_52_Re,
  output [31:0] io_out_52_Im,
  output [31:0] io_out_53_Re,
  output [31:0] io_out_53_Im,
  output [31:0] io_out_54_Re,
  output [31:0] io_out_54_Im,
  output [31:0] io_out_55_Re,
  output [31:0] io_out_55_Im,
  output [31:0] io_out_56_Re,
  output [31:0] io_out_56_Im,
  output [31:0] io_out_57_Re,
  output [31:0] io_out_57_Im,
  output [31:0] io_out_58_Re,
  output [31:0] io_out_58_Im,
  output [31:0] io_out_59_Re,
  output [31:0] io_out_59_Im,
  output [31:0] io_out_60_Re,
  output [31:0] io_out_60_Im,
  output [31:0] io_out_61_Re,
  output [31:0] io_out_61_Im,
  output [31:0] io_out_62_Re,
  output [31:0] io_out_62_Im,
  output [31:0] io_out_63_Re,
  output [31:0] io_out_63_Im,
  output [31:0] io_out_64_Re,
  output [31:0] io_out_64_Im,
  output [31:0] io_out_65_Re,
  output [31:0] io_out_65_Im,
  output [31:0] io_out_66_Re,
  output [31:0] io_out_66_Im,
  output [31:0] io_out_67_Re,
  output [31:0] io_out_67_Im,
  output [31:0] io_out_68_Re,
  output [31:0] io_out_68_Im,
  output [31:0] io_out_69_Re,
  output [31:0] io_out_69_Im,
  output [31:0] io_out_70_Re,
  output [31:0] io_out_70_Im,
  output [31:0] io_out_71_Re,
  output [31:0] io_out_71_Im,
  output [31:0] io_out_72_Re,
  output [31:0] io_out_72_Im,
  output [31:0] io_out_73_Re,
  output [31:0] io_out_73_Im,
  output [31:0] io_out_74_Re,
  output [31:0] io_out_74_Im,
  output [31:0] io_out_75_Re,
  output [31:0] io_out_75_Im,
  output [31:0] io_out_76_Re,
  output [31:0] io_out_76_Im,
  output [31:0] io_out_77_Re,
  output [31:0] io_out_77_Im,
  output [31:0] io_out_78_Re,
  output [31:0] io_out_78_Im,
  output [31:0] io_out_79_Re,
  output [31:0] io_out_79_Im,
  output [31:0] io_out_80_Re,
  output [31:0] io_out_80_Im,
  output [31:0] io_out_81_Re,
  output [31:0] io_out_81_Im,
  output [31:0] io_out_82_Re,
  output [31:0] io_out_82_Im,
  output [31:0] io_out_83_Re,
  output [31:0] io_out_83_Im,
  output [31:0] io_out_84_Re,
  output [31:0] io_out_84_Im,
  output [31:0] io_out_85_Re,
  output [31:0] io_out_85_Im,
  output [31:0] io_out_86_Re,
  output [31:0] io_out_86_Im,
  output [31:0] io_out_87_Re,
  output [31:0] io_out_87_Im,
  output [31:0] io_out_88_Re,
  output [31:0] io_out_88_Im,
  output [31:0] io_out_89_Re,
  output [31:0] io_out_89_Im,
  output [31:0] io_out_90_Re,
  output [31:0] io_out_90_Im,
  output [31:0] io_out_91_Re,
  output [31:0] io_out_91_Im,
  output [31:0] io_out_92_Re,
  output [31:0] io_out_92_Im,
  output [31:0] io_out_93_Re,
  output [31:0] io_out_93_Im,
  output [31:0] io_out_94_Re,
  output [31:0] io_out_94_Im,
  output [31:0] io_out_95_Re,
  output [31:0] io_out_95_Im
);
  assign io_out_0_Re = io_in_0_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_0_Im = io_in_0_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Re = io_in_3_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_1_Im = io_in_3_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Re = io_in_6_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_2_Im = io_in_6_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_3_Re = io_in_9_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_3_Im = io_in_9_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_4_Re = io_in_12_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_4_Im = io_in_12_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_5_Re = io_in_15_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_5_Im = io_in_15_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_6_Re = io_in_18_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_6_Im = io_in_18_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_7_Re = io_in_21_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_7_Im = io_in_21_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_8_Re = io_in_24_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_8_Im = io_in_24_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_9_Re = io_in_27_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_9_Im = io_in_27_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_10_Re = io_in_30_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_10_Im = io_in_30_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_11_Re = io_in_33_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_11_Im = io_in_33_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_12_Re = io_in_36_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_12_Im = io_in_36_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_13_Re = io_in_39_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_13_Im = io_in_39_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_14_Re = io_in_42_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_14_Im = io_in_42_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_15_Re = io_in_45_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_15_Im = io_in_45_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_16_Re = io_in_48_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_16_Im = io_in_48_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_17_Re = io_in_51_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_17_Im = io_in_51_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_18_Re = io_in_54_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_18_Im = io_in_54_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_19_Re = io_in_57_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_19_Im = io_in_57_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_20_Re = io_in_60_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_20_Im = io_in_60_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_21_Re = io_in_63_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_21_Im = io_in_63_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_22_Re = io_in_66_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_22_Im = io_in_66_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_23_Re = io_in_69_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_23_Im = io_in_69_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_24_Re = io_in_72_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_24_Im = io_in_72_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_25_Re = io_in_75_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_25_Im = io_in_75_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_26_Re = io_in_78_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_26_Im = io_in_78_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_27_Re = io_in_81_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_27_Im = io_in_81_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_28_Re = io_in_84_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_28_Im = io_in_84_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_29_Re = io_in_87_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_29_Im = io_in_87_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_30_Re = io_in_90_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_30_Im = io_in_90_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_31_Re = io_in_93_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_31_Im = io_in_93_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_32_Re = io_in_1_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_32_Im = io_in_1_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_33_Re = io_in_4_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_33_Im = io_in_4_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_34_Re = io_in_7_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_34_Im = io_in_7_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_35_Re = io_in_10_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_35_Im = io_in_10_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_36_Re = io_in_13_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_36_Im = io_in_13_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_37_Re = io_in_16_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_37_Im = io_in_16_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_38_Re = io_in_19_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_38_Im = io_in_19_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_39_Re = io_in_22_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_39_Im = io_in_22_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_40_Re = io_in_25_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_40_Im = io_in_25_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_41_Re = io_in_28_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_41_Im = io_in_28_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_42_Re = io_in_31_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_42_Im = io_in_31_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_43_Re = io_in_34_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_43_Im = io_in_34_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_44_Re = io_in_37_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_44_Im = io_in_37_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_45_Re = io_in_40_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_45_Im = io_in_40_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_46_Re = io_in_43_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_46_Im = io_in_43_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_47_Re = io_in_46_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_47_Im = io_in_46_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_48_Re = io_in_49_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_48_Im = io_in_49_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_49_Re = io_in_52_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_49_Im = io_in_52_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_50_Re = io_in_55_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_50_Im = io_in_55_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_51_Re = io_in_58_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_51_Im = io_in_58_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_52_Re = io_in_61_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_52_Im = io_in_61_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_53_Re = io_in_64_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_53_Im = io_in_64_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_54_Re = io_in_67_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_54_Im = io_in_67_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_55_Re = io_in_70_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_55_Im = io_in_70_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_56_Re = io_in_73_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_56_Im = io_in_73_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_57_Re = io_in_76_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_57_Im = io_in_76_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_58_Re = io_in_79_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_58_Im = io_in_79_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_59_Re = io_in_82_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_59_Im = io_in_82_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_60_Re = io_in_85_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_60_Im = io_in_85_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_61_Re = io_in_88_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_61_Im = io_in_88_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_62_Re = io_in_91_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_62_Im = io_in_91_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_63_Re = io_in_94_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_63_Im = io_in_94_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_64_Re = io_in_2_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_64_Im = io_in_2_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_65_Re = io_in_5_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_65_Im = io_in_5_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_66_Re = io_in_8_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_66_Im = io_in_8_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_67_Re = io_in_11_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_67_Im = io_in_11_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_68_Re = io_in_14_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_68_Im = io_in_14_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_69_Re = io_in_17_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_69_Im = io_in_17_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_70_Re = io_in_20_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_70_Im = io_in_20_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_71_Re = io_in_23_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_71_Im = io_in_23_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_72_Re = io_in_26_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_72_Im = io_in_26_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_73_Re = io_in_29_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_73_Im = io_in_29_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_74_Re = io_in_32_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_74_Im = io_in_32_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_75_Re = io_in_35_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_75_Im = io_in_35_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_76_Re = io_in_38_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_76_Im = io_in_38_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_77_Re = io_in_41_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_77_Im = io_in_41_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_78_Re = io_in_44_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_78_Im = io_in_44_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_79_Re = io_in_47_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_79_Im = io_in_47_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_80_Re = io_in_50_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_80_Im = io_in_50_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_81_Re = io_in_53_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_81_Im = io_in_53_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_82_Re = io_in_56_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_82_Im = io_in_56_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_83_Re = io_in_59_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_83_Im = io_in_59_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_84_Re = io_in_62_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_84_Im = io_in_62_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_85_Re = io_in_65_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_85_Im = io_in_65_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_86_Re = io_in_68_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_86_Im = io_in_68_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_87_Re = io_in_71_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_87_Im = io_in_71_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_88_Re = io_in_74_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_88_Im = io_in_74_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_89_Re = io_in_77_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_89_Im = io_in_77_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_90_Re = io_in_80_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_90_Im = io_in_80_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_91_Re = io_in_83_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_91_Im = io_in_83_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_92_Re = io_in_86_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_92_Im = io_in_86_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_93_Re = io_in_89_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_93_Im = io_in_89_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_94_Re = io_in_92_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_94_Im = io_in_92_Im; // @[FFTDesigns.scala 2315:17]
  assign io_out_95_Re = io_in_95_Re; // @[FFTDesigns.scala 2315:17]
  assign io_out_95_Im = io_in_95_Im; // @[FFTDesigns.scala 2315:17]
endmodule
module FPComplexMult_reducable_7(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  FP_subber_clock; // @[FPComplex.scala 162:24]
  wire  FP_subber_reset; // @[FPComplex.scala 162:24]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 162:24]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 162:24]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 162:24]
  wire  FP_adder_clock; // @[FPComplex.scala 163:24]
  wire  FP_adder_reset; // @[FPComplex.scala 163:24]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 163:24]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 163:24]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 163:24]
  wire  FP_multiplier_clock; // @[FPComplex.scala 221:28]
  wire  FP_multiplier_reset; // @[FPComplex.scala 221:28]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 221:28]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 221:28]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 221:28]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 221:28]
  wire  FP_multiplier_1_reset; // @[FPComplex.scala 221:28]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 221:28]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 221:28]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 221:28]
  wire  sign_0 = io_in_a_Re[31]; // @[FPComplex.scala 165:26]
  wire  sign_1 = io_in_a_Im[31]; // @[FPComplex.scala 166:26]
  wire [7:0] exp_0 = io_in_a_Re[30:23]; // @[FPComplex.scala 168:25]
  wire [7:0] exp_1 = io_in_a_Im[30:23]; // @[FPComplex.scala 169:25]
  wire [22:0] frac_0 = io_in_a_Re[22:0]; // @[FPComplex.scala 171:26]
  wire [22:0] frac_1 = io_in_a_Im[22:0]; // @[FPComplex.scala 172:26]
  wire  new_sign_1 = sign_0 ^ io_in_b_Im[31]; // @[FPComplex.scala 181:28]
  wire  new_sign_2 = sign_1 ^ io_in_b_Im[31]; // @[FPComplex.scala 182:28]
  wire  _T = exp_0 != 8'h0; // @[FPComplex.scala 185:19]
  wire  _T_1 = exp_1 != 8'h0; // @[FPComplex.scala 190:19]
  wire [7:0] _new_exp1_0_T_3 = exp_0 - 8'h1; // @[FPComplex.scala 197:31]
  wire [7:0] new_exp1_0 = _T ? _new_exp1_0_T_3 : exp_0; // @[FPComplex.scala 196:27 197:21 199:21]
  wire [7:0] _new_exp1_1_T_3 = exp_1 - 8'h1; // @[FPComplex.scala 202:31]
  wire [7:0] new_exp1_1 = _T_1 ? _new_exp1_1_T_3 : exp_1; // @[FPComplex.scala 201:27 202:21 204:21]
  reg [31:0] regs2_0; // @[FPComplex.scala 232:26]
  reg [31:0] regs2_1; // @[FPComplex.scala 232:26]
  wire [31:0] _regs2_0_T_1 = {new_sign_1,new_exp1_0,frac_0}; // @[FPComplex.scala 234:46]
  wire [31:0] _regs2_1_T_1 = {new_sign_2,new_exp1_1,frac_1}; // @[FPComplex.scala 235:46]
  FP_subber FP_subber ( // @[FPComplex.scala 162:24]
    .clock(FP_subber_clock),
    .reset(FP_subber_reset),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_adder FP_adder ( // @[FPComplex.scala 163:24]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 221:28]
    .clock(FP_multiplier_clock),
    .reset(FP_multiplier_reset),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 221:28]
    .clock(FP_multiplier_1_clock),
    .reset(FP_multiplier_1_reset),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 254:17]
  assign io_out_s_Im = FP_adder_io_out_s; // @[FPComplex.scala 255:17]
  assign FP_subber_clock = clock;
  assign FP_subber_reset = reset;
  assign FP_subber_io_in_a = FP_multiplier_io_out_s; // @[FPComplex.scala 211:28 228:23]
  assign FP_subber_io_in_b = regs2_1; // @[FPComplex.scala 211:28 237:23]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = regs2_0; // @[FPComplex.scala 211:28 236:23]
  assign FP_adder_io_in_b = FP_multiplier_1_io_out_s; // @[FPComplex.scala 211:28 229:23]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_reset = reset;
  assign FP_multiplier_io_in_a = io_in_a_Re; // @[FPComplex.scala 224:31]
  assign FP_multiplier_io_in_b = io_in_b_Re; // @[FPComplex.scala 225:31]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_reset = reset;
  assign FP_multiplier_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 226:31]
  assign FP_multiplier_1_io_in_b = io_in_b_Re; // @[FPComplex.scala 227:31]
  always @(posedge clock) begin
    if (reset) begin // @[FPComplex.scala 232:26]
      regs2_0 <= 32'h0; // @[FPComplex.scala 232:26]
    end else begin
      regs2_0 <= _regs2_0_T_1; // @[FPComplex.scala 234:16]
    end
    if (reset) begin // @[FPComplex.scala 232:26]
      regs2_1 <= 32'h0; // @[FPComplex.scala 232:26]
    end else begin
      regs2_1 <= _regs2_1_T_1; // @[FPComplex.scala 235:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs2_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs2_1 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMult_reducable_15(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  FP_subber_clock; // @[FPComplex.scala 162:24]
  wire  FP_subber_reset; // @[FPComplex.scala 162:24]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 162:24]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 162:24]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 162:24]
  wire  FP_adder_clock; // @[FPComplex.scala 163:24]
  wire  FP_adder_reset; // @[FPComplex.scala 163:24]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 163:24]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 163:24]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 163:24]
  wire  FP_multiplier_clock; // @[FPComplex.scala 240:28]
  wire  FP_multiplier_reset; // @[FPComplex.scala 240:28]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 240:28]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 240:28]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 240:28]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 240:28]
  wire  FP_multiplier_1_reset; // @[FPComplex.scala 240:28]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 240:28]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 240:28]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 240:28]
  wire  sign_0 = io_in_a_Re[31]; // @[FPComplex.scala 165:26]
  wire  sign_1 = io_in_a_Im[31]; // @[FPComplex.scala 166:26]
  wire [7:0] exp_0 = io_in_a_Re[30:23]; // @[FPComplex.scala 168:25]
  wire [7:0] exp_1 = io_in_a_Im[30:23]; // @[FPComplex.scala 169:25]
  wire [22:0] frac_0 = io_in_a_Re[22:0]; // @[FPComplex.scala 171:26]
  wire [22:0] frac_1 = io_in_a_Im[22:0]; // @[FPComplex.scala 172:26]
  wire  new_sign_0 = sign_0 ^ io_in_b_Re[31]; // @[FPComplex.scala 180:28]
  wire  new_sign_3 = sign_1 ^ io_in_b_Re[31]; // @[FPComplex.scala 183:28]
  wire [7:0] _new_exp1_0_T_1 = exp_0 - 8'h1; // @[FPComplex.scala 186:31]
  wire [7:0] new_exp1_0 = exp_0 != 8'h0 ? _new_exp1_0_T_1 : exp_0; // @[FPComplex.scala 185:27 186:21 188:21]
  wire [7:0] _new_exp1_1_T_1 = exp_1 - 8'h1; // @[FPComplex.scala 191:31]
  wire [7:0] new_exp1_1 = exp_1 != 8'h0 ? _new_exp1_1_T_1 : exp_1; // @[FPComplex.scala 190:27 191:21 193:21]
  reg [31:0] regs1_0; // @[FPComplex.scala 213:26]
  reg [31:0] regs1_1; // @[FPComplex.scala 213:26]
  wire [31:0] _regs1_0_T_1 = {new_sign_0,new_exp1_0,frac_0}; // @[FPComplex.scala 215:46]
  wire [31:0] _regs1_1_T_1 = {new_sign_3,new_exp1_1,frac_1}; // @[FPComplex.scala 216:46]
  FP_subber FP_subber ( // @[FPComplex.scala 162:24]
    .clock(FP_subber_clock),
    .reset(FP_subber_reset),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_adder FP_adder ( // @[FPComplex.scala 163:24]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 240:28]
    .clock(FP_multiplier_clock),
    .reset(FP_multiplier_reset),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 240:28]
    .clock(FP_multiplier_1_clock),
    .reset(FP_multiplier_1_reset),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 254:17]
  assign io_out_s_Im = FP_adder_io_out_s; // @[FPComplex.scala 255:17]
  assign FP_subber_clock = clock;
  assign FP_subber_reset = reset;
  assign FP_subber_io_in_a = regs1_0; // @[FPComplex.scala 211:28 217:23]
  assign FP_subber_io_in_b = FP_multiplier_1_io_out_s; // @[FPComplex.scala 211:28 248:23]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = FP_multiplier_io_out_s; // @[FPComplex.scala 211:28 247:23]
  assign FP_adder_io_in_b = regs1_1; // @[FPComplex.scala 211:28 218:23]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_reset = reset;
  assign FP_multiplier_io_in_a = io_in_a_Re; // @[FPComplex.scala 243:31]
  assign FP_multiplier_io_in_b = 32'hbf5db3d6; // @[FPComplex.scala 244:31]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_reset = reset;
  assign FP_multiplier_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 245:31]
  assign FP_multiplier_1_io_in_b = 32'hbf5db3d6; // @[FPComplex.scala 246:31]
  always @(posedge clock) begin
    if (reset) begin // @[FPComplex.scala 213:26]
      regs1_0 <= 32'h0; // @[FPComplex.scala 213:26]
    end else begin
      regs1_0 <= _regs1_0_T_1; // @[FPComplex.scala 215:16]
    end
    if (reset) begin // @[FPComplex.scala 213:26]
      regs1_1 <= 32'h0; // @[FPComplex.scala 213:26]
    end else begin
      regs1_1 <= _regs1_1_T_1; // @[FPComplex.scala 216:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs1_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs1_1 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactors_mr(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  input  [31:0] io_in_32_Re,
  input  [31:0] io_in_32_Im,
  input  [31:0] io_in_33_Re,
  input  [31:0] io_in_33_Im,
  input  [31:0] io_in_34_Re,
  input  [31:0] io_in_34_Im,
  input  [31:0] io_in_35_Re,
  input  [31:0] io_in_35_Im,
  input  [31:0] io_in_36_Re,
  input  [31:0] io_in_36_Im,
  input  [31:0] io_in_37_Re,
  input  [31:0] io_in_37_Im,
  input  [31:0] io_in_38_Re,
  input  [31:0] io_in_38_Im,
  input  [31:0] io_in_39_Re,
  input  [31:0] io_in_39_Im,
  input  [31:0] io_in_40_Re,
  input  [31:0] io_in_40_Im,
  input  [31:0] io_in_41_Re,
  input  [31:0] io_in_41_Im,
  input  [31:0] io_in_42_Re,
  input  [31:0] io_in_42_Im,
  input  [31:0] io_in_43_Re,
  input  [31:0] io_in_43_Im,
  input  [31:0] io_in_44_Re,
  input  [31:0] io_in_44_Im,
  input  [31:0] io_in_45_Re,
  input  [31:0] io_in_45_Im,
  input  [31:0] io_in_46_Re,
  input  [31:0] io_in_46_Im,
  input  [31:0] io_in_47_Re,
  input  [31:0] io_in_47_Im,
  input  [31:0] io_in_48_Re,
  input  [31:0] io_in_48_Im,
  input  [31:0] io_in_49_Re,
  input  [31:0] io_in_49_Im,
  input  [31:0] io_in_50_Re,
  input  [31:0] io_in_50_Im,
  input  [31:0] io_in_51_Re,
  input  [31:0] io_in_51_Im,
  input  [31:0] io_in_52_Re,
  input  [31:0] io_in_52_Im,
  input  [31:0] io_in_53_Re,
  input  [31:0] io_in_53_Im,
  input  [31:0] io_in_54_Re,
  input  [31:0] io_in_54_Im,
  input  [31:0] io_in_55_Re,
  input  [31:0] io_in_55_Im,
  input  [31:0] io_in_56_Re,
  input  [31:0] io_in_56_Im,
  input  [31:0] io_in_57_Re,
  input  [31:0] io_in_57_Im,
  input  [31:0] io_in_58_Re,
  input  [31:0] io_in_58_Im,
  input  [31:0] io_in_59_Re,
  input  [31:0] io_in_59_Im,
  input  [31:0] io_in_60_Re,
  input  [31:0] io_in_60_Im,
  input  [31:0] io_in_61_Re,
  input  [31:0] io_in_61_Im,
  input  [31:0] io_in_62_Re,
  input  [31:0] io_in_62_Im,
  input  [31:0] io_in_63_Re,
  input  [31:0] io_in_63_Im,
  input  [31:0] io_in_64_Re,
  input  [31:0] io_in_64_Im,
  input  [31:0] io_in_65_Re,
  input  [31:0] io_in_65_Im,
  input  [31:0] io_in_66_Re,
  input  [31:0] io_in_66_Im,
  input  [31:0] io_in_67_Re,
  input  [31:0] io_in_67_Im,
  input  [31:0] io_in_68_Re,
  input  [31:0] io_in_68_Im,
  input  [31:0] io_in_69_Re,
  input  [31:0] io_in_69_Im,
  input  [31:0] io_in_70_Re,
  input  [31:0] io_in_70_Im,
  input  [31:0] io_in_71_Re,
  input  [31:0] io_in_71_Im,
  input  [31:0] io_in_72_Re,
  input  [31:0] io_in_72_Im,
  input  [31:0] io_in_73_Re,
  input  [31:0] io_in_73_Im,
  input  [31:0] io_in_74_Re,
  input  [31:0] io_in_74_Im,
  input  [31:0] io_in_75_Re,
  input  [31:0] io_in_75_Im,
  input  [31:0] io_in_76_Re,
  input  [31:0] io_in_76_Im,
  input  [31:0] io_in_77_Re,
  input  [31:0] io_in_77_Im,
  input  [31:0] io_in_78_Re,
  input  [31:0] io_in_78_Im,
  input  [31:0] io_in_79_Re,
  input  [31:0] io_in_79_Im,
  input  [31:0] io_in_80_Re,
  input  [31:0] io_in_80_Im,
  input  [31:0] io_in_81_Re,
  input  [31:0] io_in_81_Im,
  input  [31:0] io_in_82_Re,
  input  [31:0] io_in_82_Im,
  input  [31:0] io_in_83_Re,
  input  [31:0] io_in_83_Im,
  input  [31:0] io_in_84_Re,
  input  [31:0] io_in_84_Im,
  input  [31:0] io_in_85_Re,
  input  [31:0] io_in_85_Im,
  input  [31:0] io_in_86_Re,
  input  [31:0] io_in_86_Im,
  input  [31:0] io_in_87_Re,
  input  [31:0] io_in_87_Im,
  input  [31:0] io_in_88_Re,
  input  [31:0] io_in_88_Im,
  input  [31:0] io_in_89_Re,
  input  [31:0] io_in_89_Im,
  input  [31:0] io_in_90_Re,
  input  [31:0] io_in_90_Im,
  input  [31:0] io_in_91_Re,
  input  [31:0] io_in_91_Im,
  input  [31:0] io_in_92_Re,
  input  [31:0] io_in_92_Im,
  input  [31:0] io_in_93_Re,
  input  [31:0] io_in_93_Im,
  input  [31:0] io_in_94_Re,
  input  [31:0] io_in_94_Im,
  input  [31:0] io_in_95_Re,
  input  [31:0] io_in_95_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im,
  output [31:0] io_out_32_Re,
  output [31:0] io_out_32_Im,
  output [31:0] io_out_33_Re,
  output [31:0] io_out_33_Im,
  output [31:0] io_out_34_Re,
  output [31:0] io_out_34_Im,
  output [31:0] io_out_35_Re,
  output [31:0] io_out_35_Im,
  output [31:0] io_out_36_Re,
  output [31:0] io_out_36_Im,
  output [31:0] io_out_37_Re,
  output [31:0] io_out_37_Im,
  output [31:0] io_out_38_Re,
  output [31:0] io_out_38_Im,
  output [31:0] io_out_39_Re,
  output [31:0] io_out_39_Im,
  output [31:0] io_out_40_Re,
  output [31:0] io_out_40_Im,
  output [31:0] io_out_41_Re,
  output [31:0] io_out_41_Im,
  output [31:0] io_out_42_Re,
  output [31:0] io_out_42_Im,
  output [31:0] io_out_43_Re,
  output [31:0] io_out_43_Im,
  output [31:0] io_out_44_Re,
  output [31:0] io_out_44_Im,
  output [31:0] io_out_45_Re,
  output [31:0] io_out_45_Im,
  output [31:0] io_out_46_Re,
  output [31:0] io_out_46_Im,
  output [31:0] io_out_47_Re,
  output [31:0] io_out_47_Im,
  output [31:0] io_out_48_Re,
  output [31:0] io_out_48_Im,
  output [31:0] io_out_49_Re,
  output [31:0] io_out_49_Im,
  output [31:0] io_out_50_Re,
  output [31:0] io_out_50_Im,
  output [31:0] io_out_51_Re,
  output [31:0] io_out_51_Im,
  output [31:0] io_out_52_Re,
  output [31:0] io_out_52_Im,
  output [31:0] io_out_53_Re,
  output [31:0] io_out_53_Im,
  output [31:0] io_out_54_Re,
  output [31:0] io_out_54_Im,
  output [31:0] io_out_55_Re,
  output [31:0] io_out_55_Im,
  output [31:0] io_out_56_Re,
  output [31:0] io_out_56_Im,
  output [31:0] io_out_57_Re,
  output [31:0] io_out_57_Im,
  output [31:0] io_out_58_Re,
  output [31:0] io_out_58_Im,
  output [31:0] io_out_59_Re,
  output [31:0] io_out_59_Im,
  output [31:0] io_out_60_Re,
  output [31:0] io_out_60_Im,
  output [31:0] io_out_61_Re,
  output [31:0] io_out_61_Im,
  output [31:0] io_out_62_Re,
  output [31:0] io_out_62_Im,
  output [31:0] io_out_63_Re,
  output [31:0] io_out_63_Im,
  output [31:0] io_out_64_Re,
  output [31:0] io_out_64_Im,
  output [31:0] io_out_65_Re,
  output [31:0] io_out_65_Im,
  output [31:0] io_out_66_Re,
  output [31:0] io_out_66_Im,
  output [31:0] io_out_67_Re,
  output [31:0] io_out_67_Im,
  output [31:0] io_out_68_Re,
  output [31:0] io_out_68_Im,
  output [31:0] io_out_69_Re,
  output [31:0] io_out_69_Im,
  output [31:0] io_out_70_Re,
  output [31:0] io_out_70_Im,
  output [31:0] io_out_71_Re,
  output [31:0] io_out_71_Im,
  output [31:0] io_out_72_Re,
  output [31:0] io_out_72_Im,
  output [31:0] io_out_73_Re,
  output [31:0] io_out_73_Im,
  output [31:0] io_out_74_Re,
  output [31:0] io_out_74_Im,
  output [31:0] io_out_75_Re,
  output [31:0] io_out_75_Im,
  output [31:0] io_out_76_Re,
  output [31:0] io_out_76_Im,
  output [31:0] io_out_77_Re,
  output [31:0] io_out_77_Im,
  output [31:0] io_out_78_Re,
  output [31:0] io_out_78_Im,
  output [31:0] io_out_79_Re,
  output [31:0] io_out_79_Im,
  output [31:0] io_out_80_Re,
  output [31:0] io_out_80_Im,
  output [31:0] io_out_81_Re,
  output [31:0] io_out_81_Im,
  output [31:0] io_out_82_Re,
  output [31:0] io_out_82_Im,
  output [31:0] io_out_83_Re,
  output [31:0] io_out_83_Im,
  output [31:0] io_out_84_Re,
  output [31:0] io_out_84_Im,
  output [31:0] io_out_85_Re,
  output [31:0] io_out_85_Im,
  output [31:0] io_out_86_Re,
  output [31:0] io_out_86_Im,
  output [31:0] io_out_87_Re,
  output [31:0] io_out_87_Im,
  output [31:0] io_out_88_Re,
  output [31:0] io_out_88_Im,
  output [31:0] io_out_89_Re,
  output [31:0] io_out_89_Im,
  output [31:0] io_out_90_Re,
  output [31:0] io_out_90_Im,
  output [31:0] io_out_91_Re,
  output [31:0] io_out_91_Im,
  output [31:0] io_out_92_Re,
  output [31:0] io_out_92_Im,
  output [31:0] io_out_93_Re,
  output [31:0] io_out_93_Im,
  output [31:0] io_out_94_Re,
  output [31:0] io_out_94_Im,
  output [31:0] io_out_95_Re,
  output [31:0] io_out_95_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] cmplx_adj_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_1_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_1_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_1_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_1_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_1_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_1_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_1_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_2_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_2_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_2_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_2_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_2_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_2_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_2_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_3_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_3_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_3_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_3_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_3_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_3_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_3_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_4_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_4_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_4_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_4_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_4_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_4_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_4_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_5_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_5_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_5_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_5_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_5_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_5_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_5_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_6_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_6_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_6_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_6_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_6_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_6_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_6_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_7_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_7_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_7_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_7_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_7_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_7_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_7_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_8_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_8_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_8_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_8_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_8_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_8_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_8_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_9_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_9_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_9_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_9_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_9_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_9_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_9_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_10_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_10_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_10_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_10_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_10_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_10_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_10_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_11_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_11_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_11_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_11_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_11_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_11_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_11_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_12_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_12_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_12_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_12_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_12_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_12_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_12_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_13_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_13_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_13_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_13_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_13_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_13_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_13_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_14_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_14_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_14_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_14_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_14_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_14_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_14_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_15_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_15_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_15_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_15_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_15_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_15_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_15_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_16_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_16_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_16_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_16_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_16_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_16_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_16_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_17_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_17_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_17_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_17_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_17_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_17_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_17_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_18_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_18_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_18_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_18_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_18_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_18_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_18_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_19_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_19_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_19_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_19_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_19_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_19_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_19_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_20_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_20_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_20_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_20_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_20_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_20_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_20_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_21_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_21_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_21_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_21_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_21_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_21_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_21_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_22_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_22_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_22_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_22_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_22_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_22_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_22_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_23_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_23_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_23_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_23_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_23_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_23_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_23_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_24_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_24_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_24_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_24_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_24_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_24_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_24_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_25_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_25_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_25_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_25_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_25_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_25_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_25_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_26_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_26_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_26_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_26_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_26_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_26_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_26_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_27_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_27_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_27_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_27_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_27_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_27_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_27_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_28_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_28_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_28_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_28_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_28_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_28_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_28_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_29_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_29_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_29_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_29_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_29_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_29_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_29_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_30_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_30_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_30_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_30_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_30_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_30_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_30_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_31_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_31_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_31_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_31_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_31_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_31_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_31_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_32_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_32_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_32_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_32_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_32_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_32_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_32_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_33_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_33_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_33_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_33_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_33_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_33_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_33_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_34_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_34_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_34_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_34_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_34_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_34_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_34_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_35_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_35_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_35_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_35_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_35_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_35_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_35_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_36_io_in_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_36_io_in_Im; // @[FFTDesigns.scala 3212:22]
  wire [7:0] cmplx_adj_36_io_in_adj; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_36_io_is_neg; // @[FFTDesigns.scala 3212:22]
  wire  cmplx_adj_36_io_is_flip; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_36_io_out_Re; // @[FFTDesigns.scala 3212:22]
  wire [31:0] cmplx_adj_36_io_out_Im; // @[FFTDesigns.scala 3212:22]
  wire  FPComplexMult_reducable_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_1_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_1_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_1_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_1_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_1_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_1_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_1_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_1_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_2_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_2_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_2_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_2_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_2_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_2_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_2_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_2_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_3_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_3_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_3_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_3_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_3_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_3_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_3_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_3_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_4_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_4_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_4_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_4_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_4_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_4_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_4_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_4_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_5_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_5_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_5_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_5_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_5_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_5_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_5_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_5_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_6_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_6_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_6_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_6_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_6_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_6_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_6_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_6_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_7_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_7_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_7_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_7_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_7_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_7_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_7_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_7_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_8_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_8_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_8_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_8_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_8_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_8_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_8_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_8_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_9_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_9_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_9_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_9_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_9_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_9_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_9_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_9_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_10_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_10_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_10_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_10_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_10_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_10_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_10_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_10_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_11_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_11_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_11_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_11_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_11_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_11_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_11_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_11_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_12_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_12_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_12_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_12_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_12_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_12_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_12_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_12_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_13_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_13_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_13_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_13_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_13_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_13_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_13_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_13_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_14_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_14_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_14_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_14_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_14_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_14_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_14_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_14_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_15_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_15_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_15_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_15_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_15_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_15_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_15_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_16_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_16_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_16_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_16_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_16_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_16_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_16_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_16_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_17_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_17_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_17_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_17_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_17_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_17_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_17_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_17_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_18_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_18_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_18_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_18_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_18_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_18_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_18_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_18_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_19_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_19_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_19_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_19_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_19_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_19_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_19_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_19_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_20_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_20_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_20_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_20_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_20_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_20_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_20_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_20_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_21_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_21_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_21_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_21_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_21_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_21_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_21_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_21_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_22_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_22_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_22_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_22_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_22_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_22_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_22_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_22_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_23_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_23_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_23_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_23_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_23_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_23_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_23_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_23_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_24_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_24_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_24_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_24_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_24_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_24_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_24_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_24_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_25_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_25_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_25_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_25_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_25_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_25_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_25_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_25_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_26_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_26_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_26_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_26_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_26_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_26_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_26_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_26_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_27_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_27_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_27_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_27_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_27_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_27_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_27_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_27_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_28_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_28_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_28_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_28_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_28_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_28_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_28_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_28_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_29_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_29_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_29_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_29_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_29_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_29_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_29_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_29_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_30_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_30_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_30_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_30_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_30_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_30_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_30_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_30_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_31_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_31_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_31_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_31_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_31_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_31_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_31_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_31_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_32_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_32_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_32_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_32_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_32_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_32_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_32_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_32_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_33_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_33_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_33_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_33_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_33_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_33_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_33_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_33_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_34_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_34_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_34_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_34_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_34_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_34_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_34_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_34_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_35_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_35_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_35_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_35_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_35_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_35_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_35_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_35_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_36_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_36_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_36_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_36_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_36_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_36_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_36_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_36_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_37_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_37_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_37_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_37_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_37_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_37_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_37_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_38_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_38_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_38_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_38_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_38_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_38_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_38_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_38_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_39_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_39_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_39_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_39_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_39_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_39_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_39_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_39_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_40_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_40_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_40_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_40_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_40_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_40_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_40_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_40_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_41_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_41_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_41_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_41_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_41_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_41_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_41_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_41_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_42_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_42_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_42_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_42_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_42_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_42_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_42_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_42_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_43_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_43_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_43_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_43_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_43_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_43_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_43_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_43_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_44_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_44_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_44_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_44_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_44_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_44_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_44_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_45_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_45_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_45_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_45_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_45_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_45_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_45_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_45_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_46_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_46_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_46_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_46_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_46_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_46_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_46_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_46_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_47_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_47_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_47_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_47_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_47_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_47_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_47_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_47_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_48_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_48_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_48_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_48_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_48_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_48_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_48_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_48_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_49_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_49_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_49_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_49_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_49_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_49_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_49_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_49_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_50_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_50_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_50_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_50_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_50_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_50_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_50_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_50_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_51_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_51_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_51_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_51_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_51_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_51_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_51_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_51_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_52_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_52_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_52_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_52_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_52_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_52_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_52_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_52_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_53_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_53_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_53_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_53_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_53_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_53_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_53_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_53_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_54_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_54_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_54_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_54_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_54_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_54_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_54_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_54_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_55_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_55_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_55_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_55_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_55_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_55_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_55_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_55_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_56_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_56_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_56_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_56_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_56_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_56_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_56_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_56_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_57_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_57_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_57_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_57_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_57_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_57_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_57_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_57_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_58_clock; // @[FFTDesigns.scala 3228:28]
  wire  FPComplexMult_reducable_58_reset; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_58_io_in_a_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_58_io_in_a_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_58_io_in_b_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_58_io_in_b_Im; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_58_io_out_s_Re; // @[FFTDesigns.scala 3228:28]
  wire [31:0] FPComplexMult_reducable_58_io_out_s_Im; // @[FFTDesigns.scala 3228:28]
  reg [31:0] reg_syncs_0_0_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_0_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_1_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_1_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_2_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_2_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_3_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_3_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_4_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_4_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_5_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_5_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_6_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_6_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_7_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_7_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_8_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_8_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_9_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_9_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_10_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_10_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_11_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_11_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_12_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_12_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_13_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_13_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_14_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_14_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_15_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_15_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_16_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_16_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_17_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_17_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_18_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_18_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_19_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_19_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_20_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_20_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_21_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_21_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_22_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_22_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_23_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_23_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_24_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_24_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_25_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_25_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_26_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_26_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_27_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_27_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_28_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_28_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_29_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_29_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_30_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_30_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_31_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_31_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_32_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_32_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_33_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_33_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_34_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_34_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_35_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_35_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_36_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_0_36_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_0_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_0_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_1_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_1_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_2_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_2_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_3_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_3_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_4_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_4_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_5_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_5_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_6_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_6_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_7_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_7_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_8_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_8_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_9_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_9_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_10_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_10_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_11_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_11_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_12_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_12_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_13_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_13_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_14_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_14_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_15_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_15_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_16_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_16_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_17_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_17_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_18_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_18_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_19_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_19_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_20_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_20_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_21_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_21_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_22_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_22_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_23_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_23_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_24_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_24_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_25_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_25_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_26_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_26_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_27_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_27_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_28_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_28_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_29_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_29_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_30_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_30_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_31_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_31_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_32_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_32_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_33_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_33_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_34_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_34_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_35_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_35_Im; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_36_Re; // @[FFTDesigns.scala 3238:27]
  reg [31:0] reg_syncs_1_36_Im; // @[FFTDesigns.scala 3238:27]
  wire [31:0] adj_wire_0_Re = cmplx_adj_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_0_Im = cmplx_adj_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_1_Re = cmplx_adj_1_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_1_Im = cmplx_adj_1_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_2_Re = cmplx_adj_2_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_2_Im = cmplx_adj_2_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_3_Re = cmplx_adj_3_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_3_Im = cmplx_adj_3_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_4_Re = cmplx_adj_4_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_4_Im = cmplx_adj_4_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_5_Re = cmplx_adj_5_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_5_Im = cmplx_adj_5_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_6_Re = cmplx_adj_6_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_6_Im = cmplx_adj_6_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_7_Re = cmplx_adj_7_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_7_Im = cmplx_adj_7_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_8_Re = cmplx_adj_8_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_8_Im = cmplx_adj_8_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_9_Re = cmplx_adj_9_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_9_Im = cmplx_adj_9_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_10_Re = cmplx_adj_10_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_10_Im = cmplx_adj_10_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_11_Re = cmplx_adj_11_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_11_Im = cmplx_adj_11_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_12_Re = cmplx_adj_12_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_12_Im = cmplx_adj_12_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_13_Re = cmplx_adj_13_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_13_Im = cmplx_adj_13_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_14_Re = cmplx_adj_14_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_14_Im = cmplx_adj_14_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_15_Re = cmplx_adj_15_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_15_Im = cmplx_adj_15_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_16_Re = cmplx_adj_16_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_16_Im = cmplx_adj_16_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_17_Re = cmplx_adj_17_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_17_Im = cmplx_adj_17_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_18_Re = cmplx_adj_18_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_18_Im = cmplx_adj_18_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_19_Re = cmplx_adj_19_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_19_Im = cmplx_adj_19_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_20_Re = cmplx_adj_20_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_20_Im = cmplx_adj_20_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_21_Re = cmplx_adj_21_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_21_Im = cmplx_adj_21_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_22_Re = cmplx_adj_22_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_22_Im = cmplx_adj_22_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_23_Re = cmplx_adj_23_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_23_Im = cmplx_adj_23_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_24_Re = cmplx_adj_24_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_24_Im = cmplx_adj_24_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_25_Re = cmplx_adj_25_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_25_Im = cmplx_adj_25_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_26_Re = cmplx_adj_26_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_26_Im = cmplx_adj_26_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_27_Re = cmplx_adj_27_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_27_Im = cmplx_adj_27_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_28_Re = cmplx_adj_28_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_28_Im = cmplx_adj_28_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_29_Re = cmplx_adj_29_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_29_Im = cmplx_adj_29_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_30_Re = cmplx_adj_30_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_30_Im = cmplx_adj_30_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_31_Re = cmplx_adj_31_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_31_Im = cmplx_adj_31_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_32_Re = cmplx_adj_32_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_32_Im = cmplx_adj_32_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_56_Re = cmplx_adj_33_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_56_Im = cmplx_adj_33_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_64_Re = cmplx_adj_34_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_64_Im = cmplx_adj_34_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_76_Re = cmplx_adj_35_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_76_Im = cmplx_adj_35_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_88_Re = cmplx_adj_36_io_out_Re; // @[FFTDesigns.scala 3215:24 3221:42]
  wire [31:0] adj_wire_88_Im = cmplx_adj_36_io_out_Im; // @[FFTDesigns.scala 3215:24 3221:42]
  cmplx_adj cmplx_adj ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  cmplx_adj cmplx_adj_1 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_1_io_in_Re),
    .io_in_Im(cmplx_adj_1_io_in_Im),
    .io_in_adj(cmplx_adj_1_io_in_adj),
    .io_is_neg(cmplx_adj_1_io_is_neg),
    .io_is_flip(cmplx_adj_1_io_is_flip),
    .io_out_Re(cmplx_adj_1_io_out_Re),
    .io_out_Im(cmplx_adj_1_io_out_Im)
  );
  cmplx_adj cmplx_adj_2 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_2_io_in_Re),
    .io_in_Im(cmplx_adj_2_io_in_Im),
    .io_in_adj(cmplx_adj_2_io_in_adj),
    .io_is_neg(cmplx_adj_2_io_is_neg),
    .io_is_flip(cmplx_adj_2_io_is_flip),
    .io_out_Re(cmplx_adj_2_io_out_Re),
    .io_out_Im(cmplx_adj_2_io_out_Im)
  );
  cmplx_adj cmplx_adj_3 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_3_io_in_Re),
    .io_in_Im(cmplx_adj_3_io_in_Im),
    .io_in_adj(cmplx_adj_3_io_in_adj),
    .io_is_neg(cmplx_adj_3_io_is_neg),
    .io_is_flip(cmplx_adj_3_io_is_flip),
    .io_out_Re(cmplx_adj_3_io_out_Re),
    .io_out_Im(cmplx_adj_3_io_out_Im)
  );
  cmplx_adj cmplx_adj_4 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_4_io_in_Re),
    .io_in_Im(cmplx_adj_4_io_in_Im),
    .io_in_adj(cmplx_adj_4_io_in_adj),
    .io_is_neg(cmplx_adj_4_io_is_neg),
    .io_is_flip(cmplx_adj_4_io_is_flip),
    .io_out_Re(cmplx_adj_4_io_out_Re),
    .io_out_Im(cmplx_adj_4_io_out_Im)
  );
  cmplx_adj cmplx_adj_5 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_5_io_in_Re),
    .io_in_Im(cmplx_adj_5_io_in_Im),
    .io_in_adj(cmplx_adj_5_io_in_adj),
    .io_is_neg(cmplx_adj_5_io_is_neg),
    .io_is_flip(cmplx_adj_5_io_is_flip),
    .io_out_Re(cmplx_adj_5_io_out_Re),
    .io_out_Im(cmplx_adj_5_io_out_Im)
  );
  cmplx_adj cmplx_adj_6 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_6_io_in_Re),
    .io_in_Im(cmplx_adj_6_io_in_Im),
    .io_in_adj(cmplx_adj_6_io_in_adj),
    .io_is_neg(cmplx_adj_6_io_is_neg),
    .io_is_flip(cmplx_adj_6_io_is_flip),
    .io_out_Re(cmplx_adj_6_io_out_Re),
    .io_out_Im(cmplx_adj_6_io_out_Im)
  );
  cmplx_adj cmplx_adj_7 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_7_io_in_Re),
    .io_in_Im(cmplx_adj_7_io_in_Im),
    .io_in_adj(cmplx_adj_7_io_in_adj),
    .io_is_neg(cmplx_adj_7_io_is_neg),
    .io_is_flip(cmplx_adj_7_io_is_flip),
    .io_out_Re(cmplx_adj_7_io_out_Re),
    .io_out_Im(cmplx_adj_7_io_out_Im)
  );
  cmplx_adj cmplx_adj_8 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_8_io_in_Re),
    .io_in_Im(cmplx_adj_8_io_in_Im),
    .io_in_adj(cmplx_adj_8_io_in_adj),
    .io_is_neg(cmplx_adj_8_io_is_neg),
    .io_is_flip(cmplx_adj_8_io_is_flip),
    .io_out_Re(cmplx_adj_8_io_out_Re),
    .io_out_Im(cmplx_adj_8_io_out_Im)
  );
  cmplx_adj cmplx_adj_9 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_9_io_in_Re),
    .io_in_Im(cmplx_adj_9_io_in_Im),
    .io_in_adj(cmplx_adj_9_io_in_adj),
    .io_is_neg(cmplx_adj_9_io_is_neg),
    .io_is_flip(cmplx_adj_9_io_is_flip),
    .io_out_Re(cmplx_adj_9_io_out_Re),
    .io_out_Im(cmplx_adj_9_io_out_Im)
  );
  cmplx_adj cmplx_adj_10 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_10_io_in_Re),
    .io_in_Im(cmplx_adj_10_io_in_Im),
    .io_in_adj(cmplx_adj_10_io_in_adj),
    .io_is_neg(cmplx_adj_10_io_is_neg),
    .io_is_flip(cmplx_adj_10_io_is_flip),
    .io_out_Re(cmplx_adj_10_io_out_Re),
    .io_out_Im(cmplx_adj_10_io_out_Im)
  );
  cmplx_adj cmplx_adj_11 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_11_io_in_Re),
    .io_in_Im(cmplx_adj_11_io_in_Im),
    .io_in_adj(cmplx_adj_11_io_in_adj),
    .io_is_neg(cmplx_adj_11_io_is_neg),
    .io_is_flip(cmplx_adj_11_io_is_flip),
    .io_out_Re(cmplx_adj_11_io_out_Re),
    .io_out_Im(cmplx_adj_11_io_out_Im)
  );
  cmplx_adj cmplx_adj_12 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_12_io_in_Re),
    .io_in_Im(cmplx_adj_12_io_in_Im),
    .io_in_adj(cmplx_adj_12_io_in_adj),
    .io_is_neg(cmplx_adj_12_io_is_neg),
    .io_is_flip(cmplx_adj_12_io_is_flip),
    .io_out_Re(cmplx_adj_12_io_out_Re),
    .io_out_Im(cmplx_adj_12_io_out_Im)
  );
  cmplx_adj cmplx_adj_13 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_13_io_in_Re),
    .io_in_Im(cmplx_adj_13_io_in_Im),
    .io_in_adj(cmplx_adj_13_io_in_adj),
    .io_is_neg(cmplx_adj_13_io_is_neg),
    .io_is_flip(cmplx_adj_13_io_is_flip),
    .io_out_Re(cmplx_adj_13_io_out_Re),
    .io_out_Im(cmplx_adj_13_io_out_Im)
  );
  cmplx_adj cmplx_adj_14 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_14_io_in_Re),
    .io_in_Im(cmplx_adj_14_io_in_Im),
    .io_in_adj(cmplx_adj_14_io_in_adj),
    .io_is_neg(cmplx_adj_14_io_is_neg),
    .io_is_flip(cmplx_adj_14_io_is_flip),
    .io_out_Re(cmplx_adj_14_io_out_Re),
    .io_out_Im(cmplx_adj_14_io_out_Im)
  );
  cmplx_adj cmplx_adj_15 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_15_io_in_Re),
    .io_in_Im(cmplx_adj_15_io_in_Im),
    .io_in_adj(cmplx_adj_15_io_in_adj),
    .io_is_neg(cmplx_adj_15_io_is_neg),
    .io_is_flip(cmplx_adj_15_io_is_flip),
    .io_out_Re(cmplx_adj_15_io_out_Re),
    .io_out_Im(cmplx_adj_15_io_out_Im)
  );
  cmplx_adj cmplx_adj_16 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_16_io_in_Re),
    .io_in_Im(cmplx_adj_16_io_in_Im),
    .io_in_adj(cmplx_adj_16_io_in_adj),
    .io_is_neg(cmplx_adj_16_io_is_neg),
    .io_is_flip(cmplx_adj_16_io_is_flip),
    .io_out_Re(cmplx_adj_16_io_out_Re),
    .io_out_Im(cmplx_adj_16_io_out_Im)
  );
  cmplx_adj cmplx_adj_17 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_17_io_in_Re),
    .io_in_Im(cmplx_adj_17_io_in_Im),
    .io_in_adj(cmplx_adj_17_io_in_adj),
    .io_is_neg(cmplx_adj_17_io_is_neg),
    .io_is_flip(cmplx_adj_17_io_is_flip),
    .io_out_Re(cmplx_adj_17_io_out_Re),
    .io_out_Im(cmplx_adj_17_io_out_Im)
  );
  cmplx_adj cmplx_adj_18 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_18_io_in_Re),
    .io_in_Im(cmplx_adj_18_io_in_Im),
    .io_in_adj(cmplx_adj_18_io_in_adj),
    .io_is_neg(cmplx_adj_18_io_is_neg),
    .io_is_flip(cmplx_adj_18_io_is_flip),
    .io_out_Re(cmplx_adj_18_io_out_Re),
    .io_out_Im(cmplx_adj_18_io_out_Im)
  );
  cmplx_adj cmplx_adj_19 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_19_io_in_Re),
    .io_in_Im(cmplx_adj_19_io_in_Im),
    .io_in_adj(cmplx_adj_19_io_in_adj),
    .io_is_neg(cmplx_adj_19_io_is_neg),
    .io_is_flip(cmplx_adj_19_io_is_flip),
    .io_out_Re(cmplx_adj_19_io_out_Re),
    .io_out_Im(cmplx_adj_19_io_out_Im)
  );
  cmplx_adj cmplx_adj_20 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_20_io_in_Re),
    .io_in_Im(cmplx_adj_20_io_in_Im),
    .io_in_adj(cmplx_adj_20_io_in_adj),
    .io_is_neg(cmplx_adj_20_io_is_neg),
    .io_is_flip(cmplx_adj_20_io_is_flip),
    .io_out_Re(cmplx_adj_20_io_out_Re),
    .io_out_Im(cmplx_adj_20_io_out_Im)
  );
  cmplx_adj cmplx_adj_21 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_21_io_in_Re),
    .io_in_Im(cmplx_adj_21_io_in_Im),
    .io_in_adj(cmplx_adj_21_io_in_adj),
    .io_is_neg(cmplx_adj_21_io_is_neg),
    .io_is_flip(cmplx_adj_21_io_is_flip),
    .io_out_Re(cmplx_adj_21_io_out_Re),
    .io_out_Im(cmplx_adj_21_io_out_Im)
  );
  cmplx_adj cmplx_adj_22 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_22_io_in_Re),
    .io_in_Im(cmplx_adj_22_io_in_Im),
    .io_in_adj(cmplx_adj_22_io_in_adj),
    .io_is_neg(cmplx_adj_22_io_is_neg),
    .io_is_flip(cmplx_adj_22_io_is_flip),
    .io_out_Re(cmplx_adj_22_io_out_Re),
    .io_out_Im(cmplx_adj_22_io_out_Im)
  );
  cmplx_adj cmplx_adj_23 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_23_io_in_Re),
    .io_in_Im(cmplx_adj_23_io_in_Im),
    .io_in_adj(cmplx_adj_23_io_in_adj),
    .io_is_neg(cmplx_adj_23_io_is_neg),
    .io_is_flip(cmplx_adj_23_io_is_flip),
    .io_out_Re(cmplx_adj_23_io_out_Re),
    .io_out_Im(cmplx_adj_23_io_out_Im)
  );
  cmplx_adj cmplx_adj_24 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_24_io_in_Re),
    .io_in_Im(cmplx_adj_24_io_in_Im),
    .io_in_adj(cmplx_adj_24_io_in_adj),
    .io_is_neg(cmplx_adj_24_io_is_neg),
    .io_is_flip(cmplx_adj_24_io_is_flip),
    .io_out_Re(cmplx_adj_24_io_out_Re),
    .io_out_Im(cmplx_adj_24_io_out_Im)
  );
  cmplx_adj cmplx_adj_25 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_25_io_in_Re),
    .io_in_Im(cmplx_adj_25_io_in_Im),
    .io_in_adj(cmplx_adj_25_io_in_adj),
    .io_is_neg(cmplx_adj_25_io_is_neg),
    .io_is_flip(cmplx_adj_25_io_is_flip),
    .io_out_Re(cmplx_adj_25_io_out_Re),
    .io_out_Im(cmplx_adj_25_io_out_Im)
  );
  cmplx_adj cmplx_adj_26 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_26_io_in_Re),
    .io_in_Im(cmplx_adj_26_io_in_Im),
    .io_in_adj(cmplx_adj_26_io_in_adj),
    .io_is_neg(cmplx_adj_26_io_is_neg),
    .io_is_flip(cmplx_adj_26_io_is_flip),
    .io_out_Re(cmplx_adj_26_io_out_Re),
    .io_out_Im(cmplx_adj_26_io_out_Im)
  );
  cmplx_adj cmplx_adj_27 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_27_io_in_Re),
    .io_in_Im(cmplx_adj_27_io_in_Im),
    .io_in_adj(cmplx_adj_27_io_in_adj),
    .io_is_neg(cmplx_adj_27_io_is_neg),
    .io_is_flip(cmplx_adj_27_io_is_flip),
    .io_out_Re(cmplx_adj_27_io_out_Re),
    .io_out_Im(cmplx_adj_27_io_out_Im)
  );
  cmplx_adj cmplx_adj_28 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_28_io_in_Re),
    .io_in_Im(cmplx_adj_28_io_in_Im),
    .io_in_adj(cmplx_adj_28_io_in_adj),
    .io_is_neg(cmplx_adj_28_io_is_neg),
    .io_is_flip(cmplx_adj_28_io_is_flip),
    .io_out_Re(cmplx_adj_28_io_out_Re),
    .io_out_Im(cmplx_adj_28_io_out_Im)
  );
  cmplx_adj cmplx_adj_29 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_29_io_in_Re),
    .io_in_Im(cmplx_adj_29_io_in_Im),
    .io_in_adj(cmplx_adj_29_io_in_adj),
    .io_is_neg(cmplx_adj_29_io_is_neg),
    .io_is_flip(cmplx_adj_29_io_is_flip),
    .io_out_Re(cmplx_adj_29_io_out_Re),
    .io_out_Im(cmplx_adj_29_io_out_Im)
  );
  cmplx_adj cmplx_adj_30 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_30_io_in_Re),
    .io_in_Im(cmplx_adj_30_io_in_Im),
    .io_in_adj(cmplx_adj_30_io_in_adj),
    .io_is_neg(cmplx_adj_30_io_is_neg),
    .io_is_flip(cmplx_adj_30_io_is_flip),
    .io_out_Re(cmplx_adj_30_io_out_Re),
    .io_out_Im(cmplx_adj_30_io_out_Im)
  );
  cmplx_adj cmplx_adj_31 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_31_io_in_Re),
    .io_in_Im(cmplx_adj_31_io_in_Im),
    .io_in_adj(cmplx_adj_31_io_in_adj),
    .io_is_neg(cmplx_adj_31_io_is_neg),
    .io_is_flip(cmplx_adj_31_io_is_flip),
    .io_out_Re(cmplx_adj_31_io_out_Re),
    .io_out_Im(cmplx_adj_31_io_out_Im)
  );
  cmplx_adj cmplx_adj_32 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_32_io_in_Re),
    .io_in_Im(cmplx_adj_32_io_in_Im),
    .io_in_adj(cmplx_adj_32_io_in_adj),
    .io_is_neg(cmplx_adj_32_io_is_neg),
    .io_is_flip(cmplx_adj_32_io_is_flip),
    .io_out_Re(cmplx_adj_32_io_out_Re),
    .io_out_Im(cmplx_adj_32_io_out_Im)
  );
  cmplx_adj cmplx_adj_33 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_33_io_in_Re),
    .io_in_Im(cmplx_adj_33_io_in_Im),
    .io_in_adj(cmplx_adj_33_io_in_adj),
    .io_is_neg(cmplx_adj_33_io_is_neg),
    .io_is_flip(cmplx_adj_33_io_is_flip),
    .io_out_Re(cmplx_adj_33_io_out_Re),
    .io_out_Im(cmplx_adj_33_io_out_Im)
  );
  cmplx_adj cmplx_adj_34 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_34_io_in_Re),
    .io_in_Im(cmplx_adj_34_io_in_Im),
    .io_in_adj(cmplx_adj_34_io_in_adj),
    .io_is_neg(cmplx_adj_34_io_is_neg),
    .io_is_flip(cmplx_adj_34_io_is_flip),
    .io_out_Re(cmplx_adj_34_io_out_Re),
    .io_out_Im(cmplx_adj_34_io_out_Im)
  );
  cmplx_adj cmplx_adj_35 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_35_io_in_Re),
    .io_in_Im(cmplx_adj_35_io_in_Im),
    .io_in_adj(cmplx_adj_35_io_in_adj),
    .io_is_neg(cmplx_adj_35_io_is_neg),
    .io_is_flip(cmplx_adj_35_io_is_flip),
    .io_out_Re(cmplx_adj_35_io_out_Re),
    .io_out_Im(cmplx_adj_35_io_out_Im)
  );
  cmplx_adj cmplx_adj_36 ( // @[FFTDesigns.scala 3212:22]
    .io_in_Re(cmplx_adj_36_io_in_Re),
    .io_in_Im(cmplx_adj_36_io_in_Im),
    .io_in_adj(cmplx_adj_36_io_in_adj),
    .io_is_neg(cmplx_adj_36_io_is_neg),
    .io_is_flip(cmplx_adj_36_io_is_flip),
    .io_out_Re(cmplx_adj_36_io_out_Re),
    .io_out_Im(cmplx_adj_36_io_out_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_clock),
    .reset(FPComplexMult_reducable_reset),
    .io_in_a_Re(FPComplexMult_reducable_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_1 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_1_clock),
    .reset(FPComplexMult_reducable_1_reset),
    .io_in_a_Re(FPComplexMult_reducable_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_1_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_2 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_2_clock),
    .reset(FPComplexMult_reducable_2_reset),
    .io_in_a_Re(FPComplexMult_reducable_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_3 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_3_clock),
    .reset(FPComplexMult_reducable_3_reset),
    .io_in_a_Re(FPComplexMult_reducable_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_3_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_4 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_4_clock),
    .reset(FPComplexMult_reducable_4_reset),
    .io_in_a_Re(FPComplexMult_reducable_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_4_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_5 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_5_clock),
    .reset(FPComplexMult_reducable_5_reset),
    .io_in_a_Re(FPComplexMult_reducable_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_5_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_6 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_6_clock),
    .reset(FPComplexMult_reducable_6_reset),
    .io_in_a_Re(FPComplexMult_reducable_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_6_io_out_s_Im)
  );
  FPComplexMult_reducable_7 FPComplexMult_reducable_7 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_7_clock),
    .reset(FPComplexMult_reducable_7_reset),
    .io_in_a_Re(FPComplexMult_reducable_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_7_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_8 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_8_clock),
    .reset(FPComplexMult_reducable_8_reset),
    .io_in_a_Re(FPComplexMult_reducable_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_8_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_9 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_9_clock),
    .reset(FPComplexMult_reducable_9_reset),
    .io_in_a_Re(FPComplexMult_reducable_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_9_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_10 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_10_clock),
    .reset(FPComplexMult_reducable_10_reset),
    .io_in_a_Re(FPComplexMult_reducable_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_10_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_11 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_11_clock),
    .reset(FPComplexMult_reducable_11_reset),
    .io_in_a_Re(FPComplexMult_reducable_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_11_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_12 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_12_clock),
    .reset(FPComplexMult_reducable_12_reset),
    .io_in_a_Re(FPComplexMult_reducable_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_12_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_13 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_13_clock),
    .reset(FPComplexMult_reducable_13_reset),
    .io_in_a_Re(FPComplexMult_reducable_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_13_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_14 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_14_clock),
    .reset(FPComplexMult_reducable_14_reset),
    .io_in_a_Re(FPComplexMult_reducable_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_14_io_out_s_Im)
  );
  FPComplexMult_reducable_15 FPComplexMult_reducable_15 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_15_clock),
    .reset(FPComplexMult_reducable_15_reset),
    .io_in_a_Re(FPComplexMult_reducable_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_15_io_in_b_Re),
    .io_out_s_Re(FPComplexMult_reducable_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_15_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_16 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_16_clock),
    .reset(FPComplexMult_reducable_16_reset),
    .io_in_a_Re(FPComplexMult_reducable_16_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_16_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_16_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_16_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_16_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_16_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_17 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_17_clock),
    .reset(FPComplexMult_reducable_17_reset),
    .io_in_a_Re(FPComplexMult_reducable_17_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_17_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_17_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_17_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_17_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_17_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_18 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_18_clock),
    .reset(FPComplexMult_reducable_18_reset),
    .io_in_a_Re(FPComplexMult_reducable_18_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_18_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_18_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_18_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_18_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_18_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_19 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_19_clock),
    .reset(FPComplexMult_reducable_19_reset),
    .io_in_a_Re(FPComplexMult_reducable_19_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_19_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_19_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_19_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_19_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_19_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_20 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_20_clock),
    .reset(FPComplexMult_reducable_20_reset),
    .io_in_a_Re(FPComplexMult_reducable_20_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_20_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_20_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_20_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_20_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_20_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_21 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_21_clock),
    .reset(FPComplexMult_reducable_21_reset),
    .io_in_a_Re(FPComplexMult_reducable_21_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_21_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_21_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_21_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_21_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_21_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_22 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_22_clock),
    .reset(FPComplexMult_reducable_22_reset),
    .io_in_a_Re(FPComplexMult_reducable_22_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_22_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_22_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_22_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_22_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_22_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_23 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_23_clock),
    .reset(FPComplexMult_reducable_23_reset),
    .io_in_a_Re(FPComplexMult_reducable_23_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_23_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_23_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_23_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_23_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_23_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_24 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_24_clock),
    .reset(FPComplexMult_reducable_24_reset),
    .io_in_a_Re(FPComplexMult_reducable_24_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_24_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_24_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_24_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_24_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_24_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_25 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_25_clock),
    .reset(FPComplexMult_reducable_25_reset),
    .io_in_a_Re(FPComplexMult_reducable_25_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_25_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_25_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_25_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_25_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_25_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_26 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_26_clock),
    .reset(FPComplexMult_reducable_26_reset),
    .io_in_a_Re(FPComplexMult_reducable_26_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_26_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_26_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_26_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_26_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_26_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_27 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_27_clock),
    .reset(FPComplexMult_reducable_27_reset),
    .io_in_a_Re(FPComplexMult_reducable_27_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_27_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_27_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_27_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_27_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_27_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_28 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_28_clock),
    .reset(FPComplexMult_reducable_28_reset),
    .io_in_a_Re(FPComplexMult_reducable_28_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_28_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_28_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_28_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_28_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_28_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_29 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_29_clock),
    .reset(FPComplexMult_reducable_29_reset),
    .io_in_a_Re(FPComplexMult_reducable_29_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_29_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_29_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_29_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_29_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_29_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_30 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_30_clock),
    .reset(FPComplexMult_reducable_30_reset),
    .io_in_a_Re(FPComplexMult_reducable_30_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_30_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_30_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_30_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_30_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_30_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_31 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_31_clock),
    .reset(FPComplexMult_reducable_31_reset),
    .io_in_a_Re(FPComplexMult_reducable_31_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_31_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_31_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_31_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_31_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_31_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_32 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_32_clock),
    .reset(FPComplexMult_reducable_32_reset),
    .io_in_a_Re(FPComplexMult_reducable_32_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_32_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_32_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_32_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_32_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_32_io_out_s_Im)
  );
  FPComplexMult_reducable_7 FPComplexMult_reducable_33 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_33_clock),
    .reset(FPComplexMult_reducable_33_reset),
    .io_in_a_Re(FPComplexMult_reducable_33_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_33_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_33_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_33_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_33_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_33_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_34 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_34_clock),
    .reset(FPComplexMult_reducable_34_reset),
    .io_in_a_Re(FPComplexMult_reducable_34_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_34_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_34_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_34_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_34_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_34_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_35 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_35_clock),
    .reset(FPComplexMult_reducable_35_reset),
    .io_in_a_Re(FPComplexMult_reducable_35_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_35_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_35_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_35_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_35_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_35_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_36 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_36_clock),
    .reset(FPComplexMult_reducable_36_reset),
    .io_in_a_Re(FPComplexMult_reducable_36_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_36_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_36_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_36_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_36_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_36_io_out_s_Im)
  );
  FPComplexMult_reducable_15 FPComplexMult_reducable_37 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_37_clock),
    .reset(FPComplexMult_reducable_37_reset),
    .io_in_a_Re(FPComplexMult_reducable_37_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_37_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_37_io_in_b_Re),
    .io_out_s_Re(FPComplexMult_reducable_37_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_37_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_38 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_38_clock),
    .reset(FPComplexMult_reducable_38_reset),
    .io_in_a_Re(FPComplexMult_reducable_38_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_38_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_38_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_38_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_38_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_38_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_39 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_39_clock),
    .reset(FPComplexMult_reducable_39_reset),
    .io_in_a_Re(FPComplexMult_reducable_39_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_39_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_39_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_39_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_39_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_39_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_40 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_40_clock),
    .reset(FPComplexMult_reducable_40_reset),
    .io_in_a_Re(FPComplexMult_reducable_40_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_40_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_40_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_40_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_40_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_40_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_41 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_41_clock),
    .reset(FPComplexMult_reducable_41_reset),
    .io_in_a_Re(FPComplexMult_reducable_41_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_41_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_41_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_41_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_41_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_41_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_42 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_42_clock),
    .reset(FPComplexMult_reducable_42_reset),
    .io_in_a_Re(FPComplexMult_reducable_42_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_42_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_42_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_42_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_42_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_42_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_43 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_43_clock),
    .reset(FPComplexMult_reducable_43_reset),
    .io_in_a_Re(FPComplexMult_reducable_43_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_43_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_43_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_43_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_43_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_43_io_out_s_Im)
  );
  FPComplexMult_reducable_15 FPComplexMult_reducable_44 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_44_clock),
    .reset(FPComplexMult_reducable_44_reset),
    .io_in_a_Re(FPComplexMult_reducable_44_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_44_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_44_io_in_b_Re),
    .io_out_s_Re(FPComplexMult_reducable_44_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_44_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_45 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_45_clock),
    .reset(FPComplexMult_reducable_45_reset),
    .io_in_a_Re(FPComplexMult_reducable_45_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_45_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_45_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_45_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_45_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_45_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_46 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_46_clock),
    .reset(FPComplexMult_reducable_46_reset),
    .io_in_a_Re(FPComplexMult_reducable_46_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_46_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_46_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_46_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_46_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_46_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_47 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_47_clock),
    .reset(FPComplexMult_reducable_47_reset),
    .io_in_a_Re(FPComplexMult_reducable_47_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_47_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_47_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_47_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_47_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_47_io_out_s_Im)
  );
  FPComplexMult_reducable_7 FPComplexMult_reducable_48 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_48_clock),
    .reset(FPComplexMult_reducable_48_reset),
    .io_in_a_Re(FPComplexMult_reducable_48_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_48_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_48_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_48_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_48_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_48_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_49 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_49_clock),
    .reset(FPComplexMult_reducable_49_reset),
    .io_in_a_Re(FPComplexMult_reducable_49_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_49_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_49_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_49_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_49_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_49_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_50 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_50_clock),
    .reset(FPComplexMult_reducable_50_reset),
    .io_in_a_Re(FPComplexMult_reducable_50_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_50_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_50_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_50_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_50_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_50_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_51 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_51_clock),
    .reset(FPComplexMult_reducable_51_reset),
    .io_in_a_Re(FPComplexMult_reducable_51_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_51_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_51_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_51_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_51_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_51_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_52 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_52_clock),
    .reset(FPComplexMult_reducable_52_reset),
    .io_in_a_Re(FPComplexMult_reducable_52_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_52_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_52_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_52_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_52_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_52_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_53 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_53_clock),
    .reset(FPComplexMult_reducable_53_reset),
    .io_in_a_Re(FPComplexMult_reducable_53_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_53_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_53_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_53_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_53_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_53_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_54 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_54_clock),
    .reset(FPComplexMult_reducable_54_reset),
    .io_in_a_Re(FPComplexMult_reducable_54_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_54_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_54_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_54_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_54_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_54_io_out_s_Im)
  );
  FPComplexMult_reducable_7 FPComplexMult_reducable_55 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_55_clock),
    .reset(FPComplexMult_reducable_55_reset),
    .io_in_a_Re(FPComplexMult_reducable_55_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_55_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_55_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_55_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_55_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_55_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_56 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_56_clock),
    .reset(FPComplexMult_reducable_56_reset),
    .io_in_a_Re(FPComplexMult_reducable_56_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_56_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_56_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_56_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_56_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_56_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_57 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_57_clock),
    .reset(FPComplexMult_reducable_57_reset),
    .io_in_a_Re(FPComplexMult_reducable_57_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_57_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_57_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_57_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_57_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_57_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_105 FPComplexMult_reducable_58 ( // @[FFTDesigns.scala 3228:28]
    .clock(FPComplexMult_reducable_58_clock),
    .reset(FPComplexMult_reducable_58_reset),
    .io_in_a_Re(FPComplexMult_reducable_58_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_58_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_reducable_58_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_reducable_58_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_reducable_58_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_58_io_out_s_Im)
  );
  assign io_out_0_Re = reg_syncs_1_0_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_0_Im = reg_syncs_1_0_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_1_Re = reg_syncs_1_1_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_1_Im = reg_syncs_1_1_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_2_Re = reg_syncs_1_2_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_2_Im = reg_syncs_1_2_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_3_Re = reg_syncs_1_3_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_3_Im = reg_syncs_1_3_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_4_Re = reg_syncs_1_4_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_4_Im = reg_syncs_1_4_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_5_Re = reg_syncs_1_5_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_5_Im = reg_syncs_1_5_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_6_Re = reg_syncs_1_6_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_6_Im = reg_syncs_1_6_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_7_Re = reg_syncs_1_7_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_7_Im = reg_syncs_1_7_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_8_Re = reg_syncs_1_8_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_8_Im = reg_syncs_1_8_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_9_Re = reg_syncs_1_9_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_9_Im = reg_syncs_1_9_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_10_Re = reg_syncs_1_10_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_10_Im = reg_syncs_1_10_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_11_Re = reg_syncs_1_11_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_11_Im = reg_syncs_1_11_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_12_Re = reg_syncs_1_12_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_12_Im = reg_syncs_1_12_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_13_Re = reg_syncs_1_13_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_13_Im = reg_syncs_1_13_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_14_Re = reg_syncs_1_14_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_14_Im = reg_syncs_1_14_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_15_Re = reg_syncs_1_15_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_15_Im = reg_syncs_1_15_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_16_Re = reg_syncs_1_16_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_16_Im = reg_syncs_1_16_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_17_Re = reg_syncs_1_17_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_17_Im = reg_syncs_1_17_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_18_Re = reg_syncs_1_18_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_18_Im = reg_syncs_1_18_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_19_Re = reg_syncs_1_19_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_19_Im = reg_syncs_1_19_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_20_Re = reg_syncs_1_20_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_20_Im = reg_syncs_1_20_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_21_Re = reg_syncs_1_21_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_21_Im = reg_syncs_1_21_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_22_Re = reg_syncs_1_22_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_22_Im = reg_syncs_1_22_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_23_Re = reg_syncs_1_23_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_23_Im = reg_syncs_1_23_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_24_Re = reg_syncs_1_24_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_24_Im = reg_syncs_1_24_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_25_Re = reg_syncs_1_25_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_25_Im = reg_syncs_1_25_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_26_Re = reg_syncs_1_26_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_26_Im = reg_syncs_1_26_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_27_Re = reg_syncs_1_27_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_27_Im = reg_syncs_1_27_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_28_Re = reg_syncs_1_28_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_28_Im = reg_syncs_1_28_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_29_Re = reg_syncs_1_29_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_29_Im = reg_syncs_1_29_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_30_Re = reg_syncs_1_30_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_30_Im = reg_syncs_1_30_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_31_Re = reg_syncs_1_31_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_31_Im = reg_syncs_1_31_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_32_Re = reg_syncs_1_32_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_32_Im = reg_syncs_1_32_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_33_Re = FPComplexMult_reducable_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_33_Im = FPComplexMult_reducable_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_34_Re = FPComplexMult_reducable_1_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_34_Im = FPComplexMult_reducable_1_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_35_Re = FPComplexMult_reducable_2_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_35_Im = FPComplexMult_reducable_2_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_36_Re = FPComplexMult_reducable_3_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_36_Im = FPComplexMult_reducable_3_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_37_Re = FPComplexMult_reducable_4_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_37_Im = FPComplexMult_reducable_4_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_38_Re = FPComplexMult_reducable_5_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_38_Im = FPComplexMult_reducable_5_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_39_Re = FPComplexMult_reducable_6_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_39_Im = FPComplexMult_reducable_6_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_40_Re = FPComplexMult_reducable_7_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_40_Im = FPComplexMult_reducable_7_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_41_Re = FPComplexMult_reducable_8_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_41_Im = FPComplexMult_reducable_8_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_42_Re = FPComplexMult_reducable_9_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_42_Im = FPComplexMult_reducable_9_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_43_Re = FPComplexMult_reducable_10_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_43_Im = FPComplexMult_reducable_10_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_44_Re = FPComplexMult_reducable_11_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_44_Im = FPComplexMult_reducable_11_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_45_Re = FPComplexMult_reducable_12_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_45_Im = FPComplexMult_reducable_12_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_46_Re = FPComplexMult_reducable_13_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_46_Im = FPComplexMult_reducable_13_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_47_Re = FPComplexMult_reducable_14_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_47_Im = FPComplexMult_reducable_14_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_48_Re = FPComplexMult_reducable_15_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_48_Im = FPComplexMult_reducable_15_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_49_Re = FPComplexMult_reducable_16_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_49_Im = FPComplexMult_reducable_16_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_50_Re = FPComplexMult_reducable_17_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_50_Im = FPComplexMult_reducable_17_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_51_Re = FPComplexMult_reducable_18_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_51_Im = FPComplexMult_reducable_18_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_52_Re = FPComplexMult_reducable_19_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_52_Im = FPComplexMult_reducable_19_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_53_Re = FPComplexMult_reducable_20_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_53_Im = FPComplexMult_reducable_20_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_54_Re = FPComplexMult_reducable_21_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_54_Im = FPComplexMult_reducable_21_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_55_Re = FPComplexMult_reducable_22_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_55_Im = FPComplexMult_reducable_22_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_56_Re = reg_syncs_1_33_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_56_Im = reg_syncs_1_33_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_57_Re = FPComplexMult_reducable_23_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_57_Im = FPComplexMult_reducable_23_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_58_Re = FPComplexMult_reducable_24_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_58_Im = FPComplexMult_reducable_24_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_59_Re = FPComplexMult_reducable_25_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_59_Im = FPComplexMult_reducable_25_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_60_Re = FPComplexMult_reducable_26_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_60_Im = FPComplexMult_reducable_26_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_61_Re = FPComplexMult_reducable_27_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_61_Im = FPComplexMult_reducable_27_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_62_Re = FPComplexMult_reducable_28_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_62_Im = FPComplexMult_reducable_28_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_63_Re = FPComplexMult_reducable_29_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_63_Im = FPComplexMult_reducable_29_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_64_Re = reg_syncs_1_34_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_64_Im = reg_syncs_1_34_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_65_Re = FPComplexMult_reducable_30_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_65_Im = FPComplexMult_reducable_30_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_66_Re = FPComplexMult_reducable_31_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_66_Im = FPComplexMult_reducable_31_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_67_Re = FPComplexMult_reducable_32_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_67_Im = FPComplexMult_reducable_32_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_68_Re = FPComplexMult_reducable_33_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_68_Im = FPComplexMult_reducable_33_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_69_Re = FPComplexMult_reducable_34_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_69_Im = FPComplexMult_reducable_34_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_70_Re = FPComplexMult_reducable_35_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_70_Im = FPComplexMult_reducable_35_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_71_Re = FPComplexMult_reducable_36_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_71_Im = FPComplexMult_reducable_36_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_72_Re = FPComplexMult_reducable_37_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_72_Im = FPComplexMult_reducable_37_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_73_Re = FPComplexMult_reducable_38_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_73_Im = FPComplexMult_reducable_38_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_74_Re = FPComplexMult_reducable_39_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_74_Im = FPComplexMult_reducable_39_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_75_Re = FPComplexMult_reducable_40_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_75_Im = FPComplexMult_reducable_40_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_76_Re = reg_syncs_1_35_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_76_Im = reg_syncs_1_35_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_77_Re = FPComplexMult_reducable_41_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_77_Im = FPComplexMult_reducable_41_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_78_Re = FPComplexMult_reducable_42_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_78_Im = FPComplexMult_reducable_42_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_79_Re = FPComplexMult_reducable_43_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_79_Im = FPComplexMult_reducable_43_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_80_Re = FPComplexMult_reducable_44_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_80_Im = FPComplexMult_reducable_44_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_81_Re = FPComplexMult_reducable_45_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_81_Im = FPComplexMult_reducable_45_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_82_Re = FPComplexMult_reducable_46_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_82_Im = FPComplexMult_reducable_46_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_83_Re = FPComplexMult_reducable_47_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_83_Im = FPComplexMult_reducable_47_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_84_Re = FPComplexMult_reducable_48_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_84_Im = FPComplexMult_reducable_48_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_85_Re = FPComplexMult_reducable_49_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_85_Im = FPComplexMult_reducable_49_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_86_Re = FPComplexMult_reducable_50_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_86_Im = FPComplexMult_reducable_50_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_87_Re = FPComplexMult_reducable_51_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_87_Im = FPComplexMult_reducable_51_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_88_Re = reg_syncs_1_36_Re; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_88_Im = reg_syncs_1_36_Im; // @[FFTDesigns.scala 3250:30 3252:42]
  assign io_out_89_Re = FPComplexMult_reducable_52_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_89_Im = FPComplexMult_reducable_52_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_90_Re = FPComplexMult_reducable_53_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_90_Im = FPComplexMult_reducable_53_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_91_Re = FPComplexMult_reducable_54_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_91_Im = FPComplexMult_reducable_54_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_92_Re = FPComplexMult_reducable_55_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_92_Im = FPComplexMult_reducable_55_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_93_Re = FPComplexMult_reducable_56_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_93_Im = FPComplexMult_reducable_56_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_94_Re = FPComplexMult_reducable_57_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_94_Im = FPComplexMult_reducable_57_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_95_Re = FPComplexMult_reducable_58_io_out_s_Re; // @[FFTDesigns.scala 3250:30 3255:33]
  assign io_out_95_Im = FPComplexMult_reducable_58_io_out_s_Im; // @[FFTDesigns.scala 3250:30 3255:33]
  assign cmplx_adj_io_in_Re = io_in_0_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_io_in_Im = io_in_0_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_1_io_in_Re = io_in_1_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_1_io_in_Im = io_in_1_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_1_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_1_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_1_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_2_io_in_Re = io_in_2_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_2_io_in_Im = io_in_2_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_2_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_2_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_2_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_3_io_in_Re = io_in_3_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_3_io_in_Im = io_in_3_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_3_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_3_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_3_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_4_io_in_Re = io_in_4_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_4_io_in_Im = io_in_4_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_4_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_4_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_4_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_5_io_in_Re = io_in_5_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_5_io_in_Im = io_in_5_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_5_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_5_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_5_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_6_io_in_Re = io_in_6_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_6_io_in_Im = io_in_6_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_6_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_6_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_6_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_7_io_in_Re = io_in_7_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_7_io_in_Im = io_in_7_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_7_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_7_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_7_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_8_io_in_Re = io_in_8_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_8_io_in_Im = io_in_8_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_8_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_8_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_8_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_9_io_in_Re = io_in_9_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_9_io_in_Im = io_in_9_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_9_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_9_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_9_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_10_io_in_Re = io_in_10_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_10_io_in_Im = io_in_10_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_10_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_10_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_10_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_11_io_in_Re = io_in_11_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_11_io_in_Im = io_in_11_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_11_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_11_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_11_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_12_io_in_Re = io_in_12_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_12_io_in_Im = io_in_12_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_12_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_12_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_12_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_13_io_in_Re = io_in_13_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_13_io_in_Im = io_in_13_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_13_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_13_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_13_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_14_io_in_Re = io_in_14_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_14_io_in_Im = io_in_14_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_14_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_14_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_14_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_15_io_in_Re = io_in_15_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_15_io_in_Im = io_in_15_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_15_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_15_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_15_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_16_io_in_Re = io_in_16_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_16_io_in_Im = io_in_16_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_16_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_16_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_16_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_17_io_in_Re = io_in_17_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_17_io_in_Im = io_in_17_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_17_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_17_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_17_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_18_io_in_Re = io_in_18_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_18_io_in_Im = io_in_18_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_18_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_18_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_18_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_19_io_in_Re = io_in_19_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_19_io_in_Im = io_in_19_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_19_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_19_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_19_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_20_io_in_Re = io_in_20_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_20_io_in_Im = io_in_20_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_20_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_20_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_20_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_21_io_in_Re = io_in_21_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_21_io_in_Im = io_in_21_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_21_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_21_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_21_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_22_io_in_Re = io_in_22_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_22_io_in_Im = io_in_22_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_22_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_22_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_22_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_23_io_in_Re = io_in_23_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_23_io_in_Im = io_in_23_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_23_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_23_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_23_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_24_io_in_Re = io_in_24_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_24_io_in_Im = io_in_24_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_24_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_24_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_24_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_25_io_in_Re = io_in_25_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_25_io_in_Im = io_in_25_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_25_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_25_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_25_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_26_io_in_Re = io_in_26_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_26_io_in_Im = io_in_26_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_26_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_26_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_26_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_27_io_in_Re = io_in_27_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_27_io_in_Im = io_in_27_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_27_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_27_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_27_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_28_io_in_Re = io_in_28_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_28_io_in_Im = io_in_28_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_28_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_28_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_28_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_29_io_in_Re = io_in_29_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_29_io_in_Im = io_in_29_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_29_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_29_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_29_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_30_io_in_Re = io_in_30_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_30_io_in_Im = io_in_30_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_30_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_30_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_30_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_31_io_in_Re = io_in_31_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_31_io_in_Im = io_in_31_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_31_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_31_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_31_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_32_io_in_Re = io_in_32_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_32_io_in_Im = io_in_32_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_32_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_32_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_32_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_33_io_in_Re = io_in_56_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_33_io_in_Im = io_in_56_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_33_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_33_io_is_neg = 1'h1; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_33_io_is_flip = 1'h1; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_34_io_in_Re = io_in_64_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_34_io_in_Im = io_in_64_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_34_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_34_io_is_neg = 1'h0; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_34_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_35_io_in_Re = io_in_76_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_35_io_in_Im = io_in_76_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_35_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_35_io_is_neg = 1'h1; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_35_io_is_flip = 1'h1; // @[FFTDesigns.scala 3220:32]
  assign cmplx_adj_36_io_in_Re = io_in_88_Re; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_36_io_in_Im = io_in_88_Im; // @[FFTDesigns.scala 3217:27]
  assign cmplx_adj_36_io_in_adj = 8'h0; // @[FFTDesigns.scala 3218:31]
  assign cmplx_adj_36_io_is_neg = 1'h1; // @[FFTDesigns.scala 3219:31]
  assign cmplx_adj_36_io_is_flip = 1'h0; // @[FFTDesigns.scala 3220:32]
  assign FPComplexMult_reducable_clock = clock;
  assign FPComplexMult_reducable_reset = reset;
  assign FPComplexMult_reducable_io_in_a_Re = io_in_33_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_io_in_a_Im = io_in_33_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_io_in_b_Re = 32'h3f7f73ae; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_io_in_b_Im = 32'hbd85f210; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_1_clock = clock;
  assign FPComplexMult_reducable_1_reset = reset;
  assign FPComplexMult_reducable_1_io_in_a_Re = io_in_34_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_1_io_in_a_Im = io_in_34_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_1_io_in_b_Re = 32'h3f7dcf54; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_1_io_in_b_Im = 32'hbe05a8a8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_2_clock = clock;
  assign FPComplexMult_reducable_2_reset = reset;
  assign FPComplexMult_reducable_2_io_in_a_Re = io_in_35_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_2_io_in_a_Im = io_in_35_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_2_io_in_b_Re = 32'h3f7b14be; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_2_io_in_b_Im = 32'hbe47c5c0; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_3_clock = clock;
  assign FPComplexMult_reducable_3_reset = reset;
  assign FPComplexMult_reducable_3_io_in_a_Re = io_in_36_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_3_io_in_a_Im = io_in_36_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_3_io_in_b_Re = 32'h3f7746ea; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_3_io_in_b_Im = 32'hbe8483ec; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_4_clock = clock;
  assign FPComplexMult_reducable_4_reset = reset;
  assign FPComplexMult_reducable_4_io_in_a_Re = io_in_37_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_4_io_in_a_Im = io_in_37_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_4_io_in_b_Re = 32'h3f726a02; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_4_io_in_b_Im = 32'hbea493b4; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_5_clock = clock;
  assign FPComplexMult_reducable_5_reset = reset;
  assign FPComplexMult_reducable_5_io_in_a_Re = io_in_38_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_5_io_in_a_Im = io_in_38_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_5_io_in_b_Re = 32'h3f6c835e; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_5_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_6_clock = clock;
  assign FPComplexMult_reducable_6_reset = reset;
  assign FPComplexMult_reducable_6_io_in_a_Re = io_in_39_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_6_io_in_a_Im = io_in_39_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_6_io_in_b_Re = 32'h3f659972; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_6_io_in_b_Im = 32'hbee273a8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_7_clock = clock;
  assign FPComplexMult_reducable_7_reset = reset;
  assign FPComplexMult_reducable_7_io_in_a_Re = io_in_40_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_7_io_in_a_Im = io_in_40_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_7_io_in_b_Re = 32'h3f5db3d6; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_7_io_in_b_Im = 32'hbefffffc; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_8_clock = clock;
  assign FPComplexMult_reducable_8_reset = reset;
  assign FPComplexMult_reducable_8_io_in_a_Re = io_in_41_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_8_io_in_a_Im = io_in_41_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_8_io_in_b_Re = 32'h3f54db30; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_8_io_in_b_Im = 32'hbf0e39d8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_9_clock = clock;
  assign FPComplexMult_reducable_9_reset = reset;
  assign FPComplexMult_reducable_9_io_in_a_Re = io_in_42_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_9_io_in_a_Im = io_in_42_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_9_io_in_b_Re = 32'h3f4b1934; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_9_io_in_b_Im = 32'hbf1bd7c8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_10_clock = clock;
  assign FPComplexMult_reducable_10_reset = reset;
  assign FPComplexMult_reducable_10_io_in_a_Re = io_in_43_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_10_io_in_a_Im = io_in_43_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_10_io_in_b_Re = 32'h3f407892; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_10_io_in_b_Im = 32'hbf28cae2; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_11_clock = clock;
  assign FPComplexMult_reducable_11_reset = reset;
  assign FPComplexMult_reducable_11_io_in_a_Re = io_in_44_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_11_io_in_a_Im = io_in_44_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_11_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_11_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_12_clock = clock;
  assign FPComplexMult_reducable_12_reset = reset;
  assign FPComplexMult_reducable_12_io_in_a_Re = io_in_45_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_12_io_in_a_Im = io_in_45_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_12_io_in_b_Re = 32'h3f28cae2; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_12_io_in_b_Im = 32'hbf407892; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_13_clock = clock;
  assign FPComplexMult_reducable_13_reset = reset;
  assign FPComplexMult_reducable_13_io_in_a_Re = io_in_46_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_13_io_in_a_Im = io_in_46_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_13_io_in_b_Re = 32'h3f1bd7c8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_13_io_in_b_Im = 32'hbf4b1934; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_14_clock = clock;
  assign FPComplexMult_reducable_14_reset = reset;
  assign FPComplexMult_reducable_14_io_in_a_Re = io_in_47_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_14_io_in_a_Im = io_in_47_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_14_io_in_b_Re = 32'h3f0e39d8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_14_io_in_b_Im = 32'hbf54db30; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_15_clock = clock;
  assign FPComplexMult_reducable_15_reset = reset;
  assign FPComplexMult_reducable_15_io_in_a_Re = io_in_48_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_15_io_in_a_Im = io_in_48_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_15_io_in_b_Re = 32'h3f000000; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_16_clock = clock;
  assign FPComplexMult_reducable_16_reset = reset;
  assign FPComplexMult_reducable_16_io_in_a_Re = io_in_49_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_16_io_in_a_Im = io_in_49_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_16_io_in_b_Re = 32'h3ee273a8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_16_io_in_b_Im = 32'hbf659972; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_17_clock = clock;
  assign FPComplexMult_reducable_17_reset = reset;
  assign FPComplexMult_reducable_17_io_in_a_Re = io_in_50_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_17_io_in_a_Im = io_in_50_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_17_io_in_b_Re = 32'h3ec3ef14; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_17_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_18_clock = clock;
  assign FPComplexMult_reducable_18_reset = reset;
  assign FPComplexMult_reducable_18_io_in_a_Re = io_in_51_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_18_io_in_a_Im = io_in_51_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_18_io_in_b_Re = 32'h3ea493b4; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_18_io_in_b_Im = 32'hbf726a02; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_19_clock = clock;
  assign FPComplexMult_reducable_19_reset = reset;
  assign FPComplexMult_reducable_19_io_in_a_Re = io_in_52_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_19_io_in_a_Im = io_in_52_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_19_io_in_b_Re = 32'h3e8483ec; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_19_io_in_b_Im = 32'hbf7746ea; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_20_clock = clock;
  assign FPComplexMult_reducable_20_reset = reset;
  assign FPComplexMult_reducable_20_io_in_a_Re = io_in_53_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_20_io_in_a_Im = io_in_53_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_20_io_in_b_Re = 32'h3e47c5c0; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_20_io_in_b_Im = 32'hbf7b14be; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_21_clock = clock;
  assign FPComplexMult_reducable_21_reset = reset;
  assign FPComplexMult_reducable_21_io_in_a_Re = io_in_54_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_21_io_in_a_Im = io_in_54_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_21_io_in_b_Re = 32'h3e05a8a8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_21_io_in_b_Im = 32'hbf7dcf54; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_22_clock = clock;
  assign FPComplexMult_reducable_22_reset = reset;
  assign FPComplexMult_reducable_22_io_in_a_Re = io_in_55_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_22_io_in_a_Im = io_in_55_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_22_io_in_b_Re = 32'h3d85f210; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_22_io_in_b_Im = 32'hbf7f73ae; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_23_clock = clock;
  assign FPComplexMult_reducable_23_reset = reset;
  assign FPComplexMult_reducable_23_io_in_a_Re = io_in_57_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_23_io_in_a_Im = io_in_57_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_23_io_in_b_Re = 32'hbd85f210; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_23_io_in_b_Im = 32'hbf7f73ae; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_24_clock = clock;
  assign FPComplexMult_reducable_24_reset = reset;
  assign FPComplexMult_reducable_24_io_in_a_Re = io_in_58_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_24_io_in_a_Im = io_in_58_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_24_io_in_b_Re = 32'hbe05a8a8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_24_io_in_b_Im = 32'hbf7dcf54; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_25_clock = clock;
  assign FPComplexMult_reducable_25_reset = reset;
  assign FPComplexMult_reducable_25_io_in_a_Re = io_in_59_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_25_io_in_a_Im = io_in_59_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_25_io_in_b_Re = 32'hbe47c5c0; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_25_io_in_b_Im = 32'hbf7b14be; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_26_clock = clock;
  assign FPComplexMult_reducable_26_reset = reset;
  assign FPComplexMult_reducable_26_io_in_a_Re = io_in_60_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_26_io_in_a_Im = io_in_60_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_26_io_in_b_Re = 32'hbe8483ec; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_26_io_in_b_Im = 32'hbf7746ea; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_27_clock = clock;
  assign FPComplexMult_reducable_27_reset = reset;
  assign FPComplexMult_reducable_27_io_in_a_Re = io_in_61_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_27_io_in_a_Im = io_in_61_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_27_io_in_b_Re = 32'hbea493b4; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_27_io_in_b_Im = 32'hbf726a02; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_28_clock = clock;
  assign FPComplexMult_reducable_28_reset = reset;
  assign FPComplexMult_reducable_28_io_in_a_Re = io_in_62_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_28_io_in_a_Im = io_in_62_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_28_io_in_b_Re = 32'hbec3ef14; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_28_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_29_clock = clock;
  assign FPComplexMult_reducable_29_reset = reset;
  assign FPComplexMult_reducable_29_io_in_a_Re = io_in_63_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_29_io_in_a_Im = io_in_63_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_29_io_in_b_Re = 32'hbee273a8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_29_io_in_b_Im = 32'hbf659972; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_30_clock = clock;
  assign FPComplexMult_reducable_30_reset = reset;
  assign FPComplexMult_reducable_30_io_in_a_Re = io_in_65_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_30_io_in_a_Im = io_in_65_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_30_io_in_b_Re = 32'h3f7dcf54; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_30_io_in_b_Im = 32'hbe05a8a8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_31_clock = clock;
  assign FPComplexMult_reducable_31_reset = reset;
  assign FPComplexMult_reducable_31_io_in_a_Re = io_in_66_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_31_io_in_a_Im = io_in_66_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_31_io_in_b_Re = 32'h3f7746ea; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_31_io_in_b_Im = 32'hbe8483ec; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_32_clock = clock;
  assign FPComplexMult_reducable_32_reset = reset;
  assign FPComplexMult_reducable_32_io_in_a_Re = io_in_67_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_32_io_in_a_Im = io_in_67_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_32_io_in_b_Re = 32'h3f6c835e; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_32_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_33_clock = clock;
  assign FPComplexMult_reducable_33_reset = reset;
  assign FPComplexMult_reducable_33_io_in_a_Re = io_in_68_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_33_io_in_a_Im = io_in_68_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_33_io_in_b_Re = 32'h3f5db3d6; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_33_io_in_b_Im = 32'hbefffffc; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_34_clock = clock;
  assign FPComplexMult_reducable_34_reset = reset;
  assign FPComplexMult_reducable_34_io_in_a_Re = io_in_69_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_34_io_in_a_Im = io_in_69_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_34_io_in_b_Re = 32'h3f4b1934; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_34_io_in_b_Im = 32'hbf1bd7c8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_35_clock = clock;
  assign FPComplexMult_reducable_35_reset = reset;
  assign FPComplexMult_reducable_35_io_in_a_Re = io_in_70_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_35_io_in_a_Im = io_in_70_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_35_io_in_b_Re = 32'h3f3504f2; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_35_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_36_clock = clock;
  assign FPComplexMult_reducable_36_reset = reset;
  assign FPComplexMult_reducable_36_io_in_a_Re = io_in_71_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_36_io_in_a_Im = io_in_71_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_36_io_in_b_Re = 32'h3f1bd7c8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_36_io_in_b_Im = 32'hbf4b1934; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_37_clock = clock;
  assign FPComplexMult_reducable_37_reset = reset;
  assign FPComplexMult_reducable_37_io_in_a_Re = io_in_72_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_37_io_in_a_Im = io_in_72_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_37_io_in_b_Re = 32'h3f000000; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_38_clock = clock;
  assign FPComplexMult_reducable_38_reset = reset;
  assign FPComplexMult_reducable_38_io_in_a_Re = io_in_73_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_38_io_in_a_Im = io_in_73_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_38_io_in_b_Re = 32'h3ec3ef14; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_38_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_39_clock = clock;
  assign FPComplexMult_reducable_39_reset = reset;
  assign FPComplexMult_reducable_39_io_in_a_Re = io_in_74_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_39_io_in_a_Im = io_in_74_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_39_io_in_b_Re = 32'h3e8483ec; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_39_io_in_b_Im = 32'hbf7746ea; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_40_clock = clock;
  assign FPComplexMult_reducable_40_reset = reset;
  assign FPComplexMult_reducable_40_io_in_a_Re = io_in_75_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_40_io_in_a_Im = io_in_75_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_40_io_in_b_Re = 32'h3e05a8a8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_40_io_in_b_Im = 32'hbf7dcf54; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_41_clock = clock;
  assign FPComplexMult_reducable_41_reset = reset;
  assign FPComplexMult_reducable_41_io_in_a_Re = io_in_77_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_41_io_in_a_Im = io_in_77_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_41_io_in_b_Re = 32'hbe05a8a8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_41_io_in_b_Im = 32'hbf7dcf54; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_42_clock = clock;
  assign FPComplexMult_reducable_42_reset = reset;
  assign FPComplexMult_reducable_42_io_in_a_Re = io_in_78_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_42_io_in_a_Im = io_in_78_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_42_io_in_b_Re = 32'hbe8483ec; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_42_io_in_b_Im = 32'hbf7746ea; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_43_clock = clock;
  assign FPComplexMult_reducable_43_reset = reset;
  assign FPComplexMult_reducable_43_io_in_a_Re = io_in_79_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_43_io_in_a_Im = io_in_79_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_43_io_in_b_Re = 32'hbec3ef14; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_43_io_in_b_Im = 32'hbf6c835e; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_44_clock = clock;
  assign FPComplexMult_reducable_44_reset = reset;
  assign FPComplexMult_reducable_44_io_in_a_Re = io_in_80_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_44_io_in_a_Im = io_in_80_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_44_io_in_b_Re = 32'hbefffffc; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_45_clock = clock;
  assign FPComplexMult_reducable_45_reset = reset;
  assign FPComplexMult_reducable_45_io_in_a_Re = io_in_81_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_45_io_in_a_Im = io_in_81_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_45_io_in_b_Re = 32'hbf1bd7c8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_45_io_in_b_Im = 32'hbf4b1934; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_46_clock = clock;
  assign FPComplexMult_reducable_46_reset = reset;
  assign FPComplexMult_reducable_46_io_in_a_Re = io_in_82_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_46_io_in_a_Im = io_in_82_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_46_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_46_io_in_b_Im = 32'hbf3504f2; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_47_clock = clock;
  assign FPComplexMult_reducable_47_reset = reset;
  assign FPComplexMult_reducable_47_io_in_a_Re = io_in_83_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_47_io_in_a_Im = io_in_83_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_47_io_in_b_Re = 32'hbf4b1934; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_47_io_in_b_Im = 32'hbf1bd7c8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_48_clock = clock;
  assign FPComplexMult_reducable_48_reset = reset;
  assign FPComplexMult_reducable_48_io_in_a_Re = io_in_84_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_48_io_in_a_Im = io_in_84_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_48_io_in_b_Re = 32'hbf5db3d6; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_48_io_in_b_Im = 32'hbf000000; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_49_clock = clock;
  assign FPComplexMult_reducable_49_reset = reset;
  assign FPComplexMult_reducable_49_io_in_a_Re = io_in_85_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_49_io_in_a_Im = io_in_85_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_49_io_in_b_Re = 32'hbf6c835e; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_49_io_in_b_Im = 32'hbec3ef14; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_50_clock = clock;
  assign FPComplexMult_reducable_50_reset = reset;
  assign FPComplexMult_reducable_50_io_in_a_Re = io_in_86_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_50_io_in_a_Im = io_in_86_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_50_io_in_b_Re = 32'hbf7746ea; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_50_io_in_b_Im = 32'hbe8483ec; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_51_clock = clock;
  assign FPComplexMult_reducable_51_reset = reset;
  assign FPComplexMult_reducable_51_io_in_a_Re = io_in_87_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_51_io_in_a_Im = io_in_87_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_51_io_in_b_Re = 32'hbf7dcf54; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_51_io_in_b_Im = 32'hbe05a8a8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_52_clock = clock;
  assign FPComplexMult_reducable_52_reset = reset;
  assign FPComplexMult_reducable_52_io_in_a_Re = io_in_89_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_52_io_in_a_Im = io_in_89_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_52_io_in_b_Re = 32'hbf7dcf54; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_52_io_in_b_Im = 32'h3e05a8a8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_53_clock = clock;
  assign FPComplexMult_reducable_53_reset = reset;
  assign FPComplexMult_reducable_53_io_in_a_Re = io_in_90_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_53_io_in_a_Im = io_in_90_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_53_io_in_b_Re = 32'hbf7746ea; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_53_io_in_b_Im = 32'h3e8483ec; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_54_clock = clock;
  assign FPComplexMult_reducable_54_reset = reset;
  assign FPComplexMult_reducable_54_io_in_a_Re = io_in_91_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_54_io_in_a_Im = io_in_91_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_54_io_in_b_Re = 32'hbf6c835e; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_54_io_in_b_Im = 32'h3ec3ef14; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_55_clock = clock;
  assign FPComplexMult_reducable_55_reset = reset;
  assign FPComplexMult_reducable_55_io_in_a_Re = io_in_92_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_55_io_in_a_Im = io_in_92_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_55_io_in_b_Re = 32'hbf5db3d6; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_55_io_in_b_Im = 32'h3efffffc; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_56_clock = clock;
  assign FPComplexMult_reducable_56_reset = reset;
  assign FPComplexMult_reducable_56_io_in_a_Re = io_in_93_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_56_io_in_a_Im = io_in_93_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_56_io_in_b_Re = 32'hbf4b1934; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_56_io_in_b_Im = 32'h3f1bd7c8; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_57_clock = clock;
  assign FPComplexMult_reducable_57_reset = reset;
  assign FPComplexMult_reducable_57_io_in_a_Re = io_in_94_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_57_io_in_a_Im = io_in_94_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_57_io_in_b_Re = 32'hbf3504f2; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_57_io_in_b_Im = 32'h3f3504f2; // @[FFTDesigns.scala 3234:28]
  assign FPComplexMult_reducable_58_clock = clock;
  assign FPComplexMult_reducable_58_reset = reset;
  assign FPComplexMult_reducable_58_io_in_a_Re = io_in_95_Re; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_58_io_in_a_Im = io_in_95_Im; // @[FFTDesigns.scala 3215:24 3224:33]
  assign FPComplexMult_reducable_58_io_in_b_Re = 32'hbf1bd7c8; // @[FFTDesigns.scala 3232:28]
  assign FPComplexMult_reducable_58_io_in_b_Im = 32'h3f4b1934; // @[FFTDesigns.scala 3234:28]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_0_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_0_Re <= adj_wire_0_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_0_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_0_Im <= adj_wire_0_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_1_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_1_Re <= adj_wire_1_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_1_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_1_Im <= adj_wire_1_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_2_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_2_Re <= adj_wire_2_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_2_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_2_Im <= adj_wire_2_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_3_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_3_Re <= adj_wire_3_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_3_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_3_Im <= adj_wire_3_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_4_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_4_Re <= adj_wire_4_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_4_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_4_Im <= adj_wire_4_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_5_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_5_Re <= adj_wire_5_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_5_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_5_Im <= adj_wire_5_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_6_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_6_Re <= adj_wire_6_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_6_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_6_Im <= adj_wire_6_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_7_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_7_Re <= adj_wire_7_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_7_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_7_Im <= adj_wire_7_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_8_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_8_Re <= adj_wire_8_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_8_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_8_Im <= adj_wire_8_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_9_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_9_Re <= adj_wire_9_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_9_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_9_Im <= adj_wire_9_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_10_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_10_Re <= adj_wire_10_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_10_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_10_Im <= adj_wire_10_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_11_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_11_Re <= adj_wire_11_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_11_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_11_Im <= adj_wire_11_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_12_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_12_Re <= adj_wire_12_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_12_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_12_Im <= adj_wire_12_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_13_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_13_Re <= adj_wire_13_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_13_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_13_Im <= adj_wire_13_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_14_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_14_Re <= adj_wire_14_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_14_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_14_Im <= adj_wire_14_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_15_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_15_Re <= adj_wire_15_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_15_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_15_Im <= adj_wire_15_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_16_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_16_Re <= adj_wire_16_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_16_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_16_Im <= adj_wire_16_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_17_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_17_Re <= adj_wire_17_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_17_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_17_Im <= adj_wire_17_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_18_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_18_Re <= adj_wire_18_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_18_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_18_Im <= adj_wire_18_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_19_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_19_Re <= adj_wire_19_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_19_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_19_Im <= adj_wire_19_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_20_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_20_Re <= adj_wire_20_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_20_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_20_Im <= adj_wire_20_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_21_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_21_Re <= adj_wire_21_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_21_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_21_Im <= adj_wire_21_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_22_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_22_Re <= adj_wire_22_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_22_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_22_Im <= adj_wire_22_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_23_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_23_Re <= adj_wire_23_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_23_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_23_Im <= adj_wire_23_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_24_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_24_Re <= adj_wire_24_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_24_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_24_Im <= adj_wire_24_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_25_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_25_Re <= adj_wire_25_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_25_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_25_Im <= adj_wire_25_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_26_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_26_Re <= adj_wire_26_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_26_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_26_Im <= adj_wire_26_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_27_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_27_Re <= adj_wire_27_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_27_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_27_Im <= adj_wire_27_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_28_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_28_Re <= adj_wire_28_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_28_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_28_Im <= adj_wire_28_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_29_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_29_Re <= adj_wire_29_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_29_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_29_Im <= adj_wire_29_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_30_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_30_Re <= adj_wire_30_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_30_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_30_Im <= adj_wire_30_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_31_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_31_Re <= adj_wire_31_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_31_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_31_Im <= adj_wire_31_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_32_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_32_Re <= adj_wire_32_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_32_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_32_Im <= adj_wire_32_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_33_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_33_Re <= adj_wire_56_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_33_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_33_Im <= adj_wire_56_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_34_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_34_Re <= adj_wire_64_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_34_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_34_Im <= adj_wire_64_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_35_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_35_Re <= adj_wire_76_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_35_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_35_Im <= adj_wire_76_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_36_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_36_Re <= adj_wire_88_Re; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_0_36_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_0_36_Im <= adj_wire_88_Im; // @[FFTDesigns.scala 3244:29]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_0_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_0_Re <= reg_syncs_0_0_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_0_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_0_Im <= reg_syncs_0_0_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_1_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_1_Re <= reg_syncs_0_1_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_1_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_1_Im <= reg_syncs_0_1_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_2_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_2_Re <= reg_syncs_0_2_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_2_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_2_Im <= reg_syncs_0_2_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_3_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_3_Re <= reg_syncs_0_3_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_3_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_3_Im <= reg_syncs_0_3_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_4_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_4_Re <= reg_syncs_0_4_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_4_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_4_Im <= reg_syncs_0_4_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_5_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_5_Re <= reg_syncs_0_5_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_5_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_5_Im <= reg_syncs_0_5_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_6_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_6_Re <= reg_syncs_0_6_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_6_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_6_Im <= reg_syncs_0_6_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_7_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_7_Re <= reg_syncs_0_7_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_7_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_7_Im <= reg_syncs_0_7_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_8_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_8_Re <= reg_syncs_0_8_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_8_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_8_Im <= reg_syncs_0_8_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_9_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_9_Re <= reg_syncs_0_9_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_9_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_9_Im <= reg_syncs_0_9_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_10_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_10_Re <= reg_syncs_0_10_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_10_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_10_Im <= reg_syncs_0_10_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_11_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_11_Re <= reg_syncs_0_11_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_11_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_11_Im <= reg_syncs_0_11_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_12_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_12_Re <= reg_syncs_0_12_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_12_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_12_Im <= reg_syncs_0_12_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_13_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_13_Re <= reg_syncs_0_13_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_13_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_13_Im <= reg_syncs_0_13_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_14_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_14_Re <= reg_syncs_0_14_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_14_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_14_Im <= reg_syncs_0_14_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_15_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_15_Re <= reg_syncs_0_15_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_15_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_15_Im <= reg_syncs_0_15_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_16_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_16_Re <= reg_syncs_0_16_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_16_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_16_Im <= reg_syncs_0_16_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_17_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_17_Re <= reg_syncs_0_17_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_17_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_17_Im <= reg_syncs_0_17_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_18_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_18_Re <= reg_syncs_0_18_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_18_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_18_Im <= reg_syncs_0_18_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_19_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_19_Re <= reg_syncs_0_19_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_19_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_19_Im <= reg_syncs_0_19_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_20_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_20_Re <= reg_syncs_0_20_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_20_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_20_Im <= reg_syncs_0_20_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_21_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_21_Re <= reg_syncs_0_21_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_21_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_21_Im <= reg_syncs_0_21_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_22_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_22_Re <= reg_syncs_0_22_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_22_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_22_Im <= reg_syncs_0_22_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_23_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_23_Re <= reg_syncs_0_23_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_23_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_23_Im <= reg_syncs_0_23_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_24_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_24_Re <= reg_syncs_0_24_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_24_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_24_Im <= reg_syncs_0_24_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_25_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_25_Re <= reg_syncs_0_25_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_25_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_25_Im <= reg_syncs_0_25_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_26_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_26_Re <= reg_syncs_0_26_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_26_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_26_Im <= reg_syncs_0_26_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_27_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_27_Re <= reg_syncs_0_27_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_27_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_27_Im <= reg_syncs_0_27_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_28_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_28_Re <= reg_syncs_0_28_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_28_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_28_Im <= reg_syncs_0_28_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_29_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_29_Re <= reg_syncs_0_29_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_29_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_29_Im <= reg_syncs_0_29_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_30_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_30_Re <= reg_syncs_0_30_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_30_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_30_Im <= reg_syncs_0_30_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_31_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_31_Re <= reg_syncs_0_31_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_31_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_31_Im <= reg_syncs_0_31_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_32_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_32_Re <= reg_syncs_0_32_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_32_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_32_Im <= reg_syncs_0_32_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_33_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_33_Re <= reg_syncs_0_33_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_33_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_33_Im <= reg_syncs_0_33_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_34_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_34_Re <= reg_syncs_0_34_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_34_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_34_Im <= reg_syncs_0_34_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_35_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_35_Re <= reg_syncs_0_35_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_35_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_35_Im <= reg_syncs_0_35_Im; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_36_Re <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_36_Re <= reg_syncs_0_36_Re; // @[FFTDesigns.scala 3247:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3238:27]
      reg_syncs_1_36_Im <= 32'h0; // @[FFTDesigns.scala 3238:27]
    end else begin
      reg_syncs_1_36_Im <= reg_syncs_0_36_Im; // @[FFTDesigns.scala 3247:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_syncs_0_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_syncs_0_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_syncs_0_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_syncs_0_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_syncs_0_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_syncs_0_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_syncs_0_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_syncs_0_3_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_syncs_0_4_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_syncs_0_4_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_syncs_0_5_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_syncs_0_5_Im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_syncs_0_6_Re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_syncs_0_6_Im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_syncs_0_7_Re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_syncs_0_7_Im = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_syncs_0_8_Re = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_syncs_0_8_Im = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_syncs_0_9_Re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_syncs_0_9_Im = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_syncs_0_10_Re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_syncs_0_10_Im = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_syncs_0_11_Re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_syncs_0_11_Im = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_syncs_0_12_Re = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_syncs_0_12_Im = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_syncs_0_13_Re = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_syncs_0_13_Im = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_syncs_0_14_Re = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_syncs_0_14_Im = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_syncs_0_15_Re = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_syncs_0_15_Im = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  reg_syncs_0_16_Re = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  reg_syncs_0_16_Im = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  reg_syncs_0_17_Re = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  reg_syncs_0_17_Im = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  reg_syncs_0_18_Re = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  reg_syncs_0_18_Im = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  reg_syncs_0_19_Re = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  reg_syncs_0_19_Im = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  reg_syncs_0_20_Re = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  reg_syncs_0_20_Im = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  reg_syncs_0_21_Re = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  reg_syncs_0_21_Im = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  reg_syncs_0_22_Re = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  reg_syncs_0_22_Im = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  reg_syncs_0_23_Re = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  reg_syncs_0_23_Im = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  reg_syncs_0_24_Re = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  reg_syncs_0_24_Im = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  reg_syncs_0_25_Re = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  reg_syncs_0_25_Im = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  reg_syncs_0_26_Re = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  reg_syncs_0_26_Im = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  reg_syncs_0_27_Re = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  reg_syncs_0_27_Im = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  reg_syncs_0_28_Re = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  reg_syncs_0_28_Im = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  reg_syncs_0_29_Re = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  reg_syncs_0_29_Im = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  reg_syncs_0_30_Re = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  reg_syncs_0_30_Im = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  reg_syncs_0_31_Re = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  reg_syncs_0_31_Im = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  reg_syncs_0_32_Re = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  reg_syncs_0_32_Im = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  reg_syncs_0_33_Re = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  reg_syncs_0_33_Im = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  reg_syncs_0_34_Re = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  reg_syncs_0_34_Im = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  reg_syncs_0_35_Re = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  reg_syncs_0_35_Im = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  reg_syncs_0_36_Re = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  reg_syncs_0_36_Im = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  reg_syncs_1_0_Re = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  reg_syncs_1_0_Im = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  reg_syncs_1_1_Re = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  reg_syncs_1_1_Im = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  reg_syncs_1_2_Re = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  reg_syncs_1_2_Im = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  reg_syncs_1_3_Re = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  reg_syncs_1_3_Im = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  reg_syncs_1_4_Re = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  reg_syncs_1_4_Im = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  reg_syncs_1_5_Re = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  reg_syncs_1_5_Im = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  reg_syncs_1_6_Re = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  reg_syncs_1_6_Im = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  reg_syncs_1_7_Re = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  reg_syncs_1_7_Im = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  reg_syncs_1_8_Re = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  reg_syncs_1_8_Im = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  reg_syncs_1_9_Re = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  reg_syncs_1_9_Im = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  reg_syncs_1_10_Re = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  reg_syncs_1_10_Im = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  reg_syncs_1_11_Re = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  reg_syncs_1_11_Im = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  reg_syncs_1_12_Re = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  reg_syncs_1_12_Im = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  reg_syncs_1_13_Re = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  reg_syncs_1_13_Im = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  reg_syncs_1_14_Re = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  reg_syncs_1_14_Im = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  reg_syncs_1_15_Re = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  reg_syncs_1_15_Im = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  reg_syncs_1_16_Re = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  reg_syncs_1_16_Im = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  reg_syncs_1_17_Re = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  reg_syncs_1_17_Im = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  reg_syncs_1_18_Re = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  reg_syncs_1_18_Im = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  reg_syncs_1_19_Re = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  reg_syncs_1_19_Im = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  reg_syncs_1_20_Re = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  reg_syncs_1_20_Im = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  reg_syncs_1_21_Re = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  reg_syncs_1_21_Im = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  reg_syncs_1_22_Re = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  reg_syncs_1_22_Im = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  reg_syncs_1_23_Re = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  reg_syncs_1_23_Im = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  reg_syncs_1_24_Re = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  reg_syncs_1_24_Im = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  reg_syncs_1_25_Re = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  reg_syncs_1_25_Im = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  reg_syncs_1_26_Re = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  reg_syncs_1_26_Im = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  reg_syncs_1_27_Re = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  reg_syncs_1_27_Im = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  reg_syncs_1_28_Re = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  reg_syncs_1_28_Im = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  reg_syncs_1_29_Re = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  reg_syncs_1_29_Im = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  reg_syncs_1_30_Re = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  reg_syncs_1_30_Im = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  reg_syncs_1_31_Re = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  reg_syncs_1_31_Im = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  reg_syncs_1_32_Re = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  reg_syncs_1_32_Im = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  reg_syncs_1_33_Re = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  reg_syncs_1_33_Im = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  reg_syncs_1_34_Re = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  reg_syncs_1_34_Im = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  reg_syncs_1_35_Re = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  reg_syncs_1_35_Im = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  reg_syncs_1_36_Re = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  reg_syncs_1_36_Im = _RAND_147[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FFT_mr96_basic(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [31:0] io_in_24_Re,
  input  [31:0] io_in_24_Im,
  input  [31:0] io_in_25_Re,
  input  [31:0] io_in_25_Im,
  input  [31:0] io_in_26_Re,
  input  [31:0] io_in_26_Im,
  input  [31:0] io_in_27_Re,
  input  [31:0] io_in_27_Im,
  input  [31:0] io_in_28_Re,
  input  [31:0] io_in_28_Im,
  input  [31:0] io_in_29_Re,
  input  [31:0] io_in_29_Im,
  input  [31:0] io_in_30_Re,
  input  [31:0] io_in_30_Im,
  input  [31:0] io_in_31_Re,
  input  [31:0] io_in_31_Im,
  input  [31:0] io_in_32_Re,
  input  [31:0] io_in_32_Im,
  input  [31:0] io_in_33_Re,
  input  [31:0] io_in_33_Im,
  input  [31:0] io_in_34_Re,
  input  [31:0] io_in_34_Im,
  input  [31:0] io_in_35_Re,
  input  [31:0] io_in_35_Im,
  input  [31:0] io_in_36_Re,
  input  [31:0] io_in_36_Im,
  input  [31:0] io_in_37_Re,
  input  [31:0] io_in_37_Im,
  input  [31:0] io_in_38_Re,
  input  [31:0] io_in_38_Im,
  input  [31:0] io_in_39_Re,
  input  [31:0] io_in_39_Im,
  input  [31:0] io_in_40_Re,
  input  [31:0] io_in_40_Im,
  input  [31:0] io_in_41_Re,
  input  [31:0] io_in_41_Im,
  input  [31:0] io_in_42_Re,
  input  [31:0] io_in_42_Im,
  input  [31:0] io_in_43_Re,
  input  [31:0] io_in_43_Im,
  input  [31:0] io_in_44_Re,
  input  [31:0] io_in_44_Im,
  input  [31:0] io_in_45_Re,
  input  [31:0] io_in_45_Im,
  input  [31:0] io_in_46_Re,
  input  [31:0] io_in_46_Im,
  input  [31:0] io_in_47_Re,
  input  [31:0] io_in_47_Im,
  input  [31:0] io_in_48_Re,
  input  [31:0] io_in_48_Im,
  input  [31:0] io_in_49_Re,
  input  [31:0] io_in_49_Im,
  input  [31:0] io_in_50_Re,
  input  [31:0] io_in_50_Im,
  input  [31:0] io_in_51_Re,
  input  [31:0] io_in_51_Im,
  input  [31:0] io_in_52_Re,
  input  [31:0] io_in_52_Im,
  input  [31:0] io_in_53_Re,
  input  [31:0] io_in_53_Im,
  input  [31:0] io_in_54_Re,
  input  [31:0] io_in_54_Im,
  input  [31:0] io_in_55_Re,
  input  [31:0] io_in_55_Im,
  input  [31:0] io_in_56_Re,
  input  [31:0] io_in_56_Im,
  input  [31:0] io_in_57_Re,
  input  [31:0] io_in_57_Im,
  input  [31:0] io_in_58_Re,
  input  [31:0] io_in_58_Im,
  input  [31:0] io_in_59_Re,
  input  [31:0] io_in_59_Im,
  input  [31:0] io_in_60_Re,
  input  [31:0] io_in_60_Im,
  input  [31:0] io_in_61_Re,
  input  [31:0] io_in_61_Im,
  input  [31:0] io_in_62_Re,
  input  [31:0] io_in_62_Im,
  input  [31:0] io_in_63_Re,
  input  [31:0] io_in_63_Im,
  input  [31:0] io_in_64_Re,
  input  [31:0] io_in_64_Im,
  input  [31:0] io_in_65_Re,
  input  [31:0] io_in_65_Im,
  input  [31:0] io_in_66_Re,
  input  [31:0] io_in_66_Im,
  input  [31:0] io_in_67_Re,
  input  [31:0] io_in_67_Im,
  input  [31:0] io_in_68_Re,
  input  [31:0] io_in_68_Im,
  input  [31:0] io_in_69_Re,
  input  [31:0] io_in_69_Im,
  input  [31:0] io_in_70_Re,
  input  [31:0] io_in_70_Im,
  input  [31:0] io_in_71_Re,
  input  [31:0] io_in_71_Im,
  input  [31:0] io_in_72_Re,
  input  [31:0] io_in_72_Im,
  input  [31:0] io_in_73_Re,
  input  [31:0] io_in_73_Im,
  input  [31:0] io_in_74_Re,
  input  [31:0] io_in_74_Im,
  input  [31:0] io_in_75_Re,
  input  [31:0] io_in_75_Im,
  input  [31:0] io_in_76_Re,
  input  [31:0] io_in_76_Im,
  input  [31:0] io_in_77_Re,
  input  [31:0] io_in_77_Im,
  input  [31:0] io_in_78_Re,
  input  [31:0] io_in_78_Im,
  input  [31:0] io_in_79_Re,
  input  [31:0] io_in_79_Im,
  input  [31:0] io_in_80_Re,
  input  [31:0] io_in_80_Im,
  input  [31:0] io_in_81_Re,
  input  [31:0] io_in_81_Im,
  input  [31:0] io_in_82_Re,
  input  [31:0] io_in_82_Im,
  input  [31:0] io_in_83_Re,
  input  [31:0] io_in_83_Im,
  input  [31:0] io_in_84_Re,
  input  [31:0] io_in_84_Im,
  input  [31:0] io_in_85_Re,
  input  [31:0] io_in_85_Im,
  input  [31:0] io_in_86_Re,
  input  [31:0] io_in_86_Im,
  input  [31:0] io_in_87_Re,
  input  [31:0] io_in_87_Im,
  input  [31:0] io_in_88_Re,
  input  [31:0] io_in_88_Im,
  input  [31:0] io_in_89_Re,
  input  [31:0] io_in_89_Im,
  input  [31:0] io_in_90_Re,
  input  [31:0] io_in_90_Im,
  input  [31:0] io_in_91_Re,
  input  [31:0] io_in_91_Im,
  input  [31:0] io_in_92_Re,
  input  [31:0] io_in_92_Im,
  input  [31:0] io_in_93_Re,
  input  [31:0] io_in_93_Im,
  input  [31:0] io_in_94_Re,
  input  [31:0] io_in_94_Im,
  input  [31:0] io_in_95_Re,
  input  [31:0] io_in_95_Im,
  input         io_in_ready,
  output        io_out_validate,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im,
  output [31:0] io_out_24_Re,
  output [31:0] io_out_24_Im,
  output [31:0] io_out_25_Re,
  output [31:0] io_out_25_Im,
  output [31:0] io_out_26_Re,
  output [31:0] io_out_26_Im,
  output [31:0] io_out_27_Re,
  output [31:0] io_out_27_Im,
  output [31:0] io_out_28_Re,
  output [31:0] io_out_28_Im,
  output [31:0] io_out_29_Re,
  output [31:0] io_out_29_Im,
  output [31:0] io_out_30_Re,
  output [31:0] io_out_30_Im,
  output [31:0] io_out_31_Re,
  output [31:0] io_out_31_Im,
  output [31:0] io_out_32_Re,
  output [31:0] io_out_32_Im,
  output [31:0] io_out_33_Re,
  output [31:0] io_out_33_Im,
  output [31:0] io_out_34_Re,
  output [31:0] io_out_34_Im,
  output [31:0] io_out_35_Re,
  output [31:0] io_out_35_Im,
  output [31:0] io_out_36_Re,
  output [31:0] io_out_36_Im,
  output [31:0] io_out_37_Re,
  output [31:0] io_out_37_Im,
  output [31:0] io_out_38_Re,
  output [31:0] io_out_38_Im,
  output [31:0] io_out_39_Re,
  output [31:0] io_out_39_Im,
  output [31:0] io_out_40_Re,
  output [31:0] io_out_40_Im,
  output [31:0] io_out_41_Re,
  output [31:0] io_out_41_Im,
  output [31:0] io_out_42_Re,
  output [31:0] io_out_42_Im,
  output [31:0] io_out_43_Re,
  output [31:0] io_out_43_Im,
  output [31:0] io_out_44_Re,
  output [31:0] io_out_44_Im,
  output [31:0] io_out_45_Re,
  output [31:0] io_out_45_Im,
  output [31:0] io_out_46_Re,
  output [31:0] io_out_46_Im,
  output [31:0] io_out_47_Re,
  output [31:0] io_out_47_Im,
  output [31:0] io_out_48_Re,
  output [31:0] io_out_48_Im,
  output [31:0] io_out_49_Re,
  output [31:0] io_out_49_Im,
  output [31:0] io_out_50_Re,
  output [31:0] io_out_50_Im,
  output [31:0] io_out_51_Re,
  output [31:0] io_out_51_Im,
  output [31:0] io_out_52_Re,
  output [31:0] io_out_52_Im,
  output [31:0] io_out_53_Re,
  output [31:0] io_out_53_Im,
  output [31:0] io_out_54_Re,
  output [31:0] io_out_54_Im,
  output [31:0] io_out_55_Re,
  output [31:0] io_out_55_Im,
  output [31:0] io_out_56_Re,
  output [31:0] io_out_56_Im,
  output [31:0] io_out_57_Re,
  output [31:0] io_out_57_Im,
  output [31:0] io_out_58_Re,
  output [31:0] io_out_58_Im,
  output [31:0] io_out_59_Re,
  output [31:0] io_out_59_Im,
  output [31:0] io_out_60_Re,
  output [31:0] io_out_60_Im,
  output [31:0] io_out_61_Re,
  output [31:0] io_out_61_Im,
  output [31:0] io_out_62_Re,
  output [31:0] io_out_62_Im,
  output [31:0] io_out_63_Re,
  output [31:0] io_out_63_Im,
  output [31:0] io_out_64_Re,
  output [31:0] io_out_64_Im,
  output [31:0] io_out_65_Re,
  output [31:0] io_out_65_Im,
  output [31:0] io_out_66_Re,
  output [31:0] io_out_66_Im,
  output [31:0] io_out_67_Re,
  output [31:0] io_out_67_Im,
  output [31:0] io_out_68_Re,
  output [31:0] io_out_68_Im,
  output [31:0] io_out_69_Re,
  output [31:0] io_out_69_Im,
  output [31:0] io_out_70_Re,
  output [31:0] io_out_70_Im,
  output [31:0] io_out_71_Re,
  output [31:0] io_out_71_Im,
  output [31:0] io_out_72_Re,
  output [31:0] io_out_72_Im,
  output [31:0] io_out_73_Re,
  output [31:0] io_out_73_Im,
  output [31:0] io_out_74_Re,
  output [31:0] io_out_74_Im,
  output [31:0] io_out_75_Re,
  output [31:0] io_out_75_Im,
  output [31:0] io_out_76_Re,
  output [31:0] io_out_76_Im,
  output [31:0] io_out_77_Re,
  output [31:0] io_out_77_Im,
  output [31:0] io_out_78_Re,
  output [31:0] io_out_78_Im,
  output [31:0] io_out_79_Re,
  output [31:0] io_out_79_Im,
  output [31:0] io_out_80_Re,
  output [31:0] io_out_80_Im,
  output [31:0] io_out_81_Re,
  output [31:0] io_out_81_Im,
  output [31:0] io_out_82_Re,
  output [31:0] io_out_82_Im,
  output [31:0] io_out_83_Re,
  output [31:0] io_out_83_Im,
  output [31:0] io_out_84_Re,
  output [31:0] io_out_84_Im,
  output [31:0] io_out_85_Re,
  output [31:0] io_out_85_Im,
  output [31:0] io_out_86_Re,
  output [31:0] io_out_86_Im,
  output [31:0] io_out_87_Re,
  output [31:0] io_out_87_Im,
  output [31:0] io_out_88_Re,
  output [31:0] io_out_88_Im,
  output [31:0] io_out_89_Re,
  output [31:0] io_out_89_Im,
  output [31:0] io_out_90_Re,
  output [31:0] io_out_90_Im,
  output [31:0] io_out_91_Re,
  output [31:0] io_out_91_Im,
  output [31:0] io_out_92_Re,
  output [31:0] io_out_92_Im,
  output [31:0] io_out_93_Re,
  output [31:0] io_out_93_Im,
  output [31:0] io_out_94_Re,
  output [31:0] io_out_94_Im,
  output [31:0] io_out_95_Re,
  output [31:0] io_out_95_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
`endif // RANDOMIZE_REG_INIT
  wire  FFT_sr_v2_nrv_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_1_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_1_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_1_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_2_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_2_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_2_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_3_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_3_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_3_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_4_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_4_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_4_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_5_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_5_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_5_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_6_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_6_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_6_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_7_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_7_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_7_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_8_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_8_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_8_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_9_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_9_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_9_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_10_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_10_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_10_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_11_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_11_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_11_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_12_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_12_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_12_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_13_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_13_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_13_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_14_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_14_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_14_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_15_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_15_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_15_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_16_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_16_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_16_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_17_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_17_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_17_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_18_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_18_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_18_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_19_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_19_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_19_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_20_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_20_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_20_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_21_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_21_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_21_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_22_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_22_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_22_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_23_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_23_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_23_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_24_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_24_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_24_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_25_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_25_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_25_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_26_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_26_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_26_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_27_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_27_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_27_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_28_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_28_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_28_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_29_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_29_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_29_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_30_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_30_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_30_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_31_clock; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_31_reset; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_in_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_in_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_in_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_in_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_in_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_in_2_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_out_0_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_out_0_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_out_1_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_out_1_Im; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_out_2_Re; // @[FFTDesigns.scala 3438:28]
  wire [31:0] FFT_sr_v2_nrv_31_io_out_2_Im; // @[FFTDesigns.scala 3438:28]
  wire  FFT_sr_v2_nrv_32_clock; // @[FFTDesigns.scala 3442:28]
  wire  FFT_sr_v2_nrv_32_reset; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_0_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_0_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_1_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_1_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_2_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_2_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_3_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_3_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_4_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_4_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_5_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_5_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_6_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_6_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_7_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_7_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_8_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_8_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_9_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_9_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_10_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_10_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_11_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_11_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_12_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_12_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_13_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_13_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_14_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_14_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_15_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_15_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_16_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_16_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_17_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_17_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_18_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_18_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_19_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_19_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_20_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_20_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_21_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_21_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_22_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_22_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_23_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_23_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_24_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_24_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_25_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_25_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_26_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_26_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_27_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_27_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_28_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_28_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_29_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_29_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_30_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_30_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_31_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_in_31_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_0_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_0_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_1_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_1_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_2_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_2_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_3_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_3_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_4_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_4_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_5_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_5_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_6_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_6_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_7_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_7_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_8_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_8_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_9_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_9_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_10_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_10_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_11_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_11_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_12_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_12_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_13_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_13_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_14_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_14_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_15_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_15_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_16_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_16_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_17_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_17_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_18_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_18_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_19_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_19_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_20_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_20_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_21_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_21_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_22_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_22_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_23_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_23_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_24_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_24_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_25_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_25_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_26_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_26_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_27_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_27_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_28_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_28_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_29_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_29_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_30_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_30_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_31_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_32_io_out_31_Im; // @[FFTDesigns.scala 3442:28]
  wire  FFT_sr_v2_nrv_33_clock; // @[FFTDesigns.scala 3442:28]
  wire  FFT_sr_v2_nrv_33_reset; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_0_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_0_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_1_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_1_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_2_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_2_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_3_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_3_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_4_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_4_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_5_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_5_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_6_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_6_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_7_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_7_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_8_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_8_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_9_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_9_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_10_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_10_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_11_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_11_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_12_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_12_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_13_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_13_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_14_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_14_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_15_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_15_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_16_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_16_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_17_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_17_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_18_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_18_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_19_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_19_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_20_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_20_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_21_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_21_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_22_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_22_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_23_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_23_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_24_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_24_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_25_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_25_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_26_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_26_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_27_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_27_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_28_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_28_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_29_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_29_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_30_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_30_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_31_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_in_31_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_0_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_0_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_1_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_1_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_2_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_2_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_3_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_3_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_4_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_4_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_5_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_5_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_6_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_6_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_7_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_7_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_8_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_8_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_9_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_9_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_10_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_10_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_11_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_11_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_12_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_12_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_13_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_13_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_14_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_14_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_15_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_15_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_16_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_16_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_17_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_17_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_18_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_18_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_19_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_19_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_20_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_20_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_21_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_21_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_22_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_22_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_23_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_23_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_24_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_24_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_25_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_25_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_26_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_26_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_27_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_27_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_28_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_28_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_29_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_29_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_30_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_30_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_31_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_33_io_out_31_Im; // @[FFTDesigns.scala 3442:28]
  wire  FFT_sr_v2_nrv_34_clock; // @[FFTDesigns.scala 3442:28]
  wire  FFT_sr_v2_nrv_34_reset; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_0_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_0_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_1_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_1_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_2_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_2_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_3_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_3_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_4_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_4_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_5_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_5_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_6_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_6_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_7_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_7_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_8_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_8_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_9_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_9_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_10_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_10_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_11_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_11_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_12_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_12_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_13_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_13_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_14_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_14_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_15_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_15_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_16_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_16_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_17_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_17_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_18_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_18_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_19_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_19_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_20_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_20_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_21_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_21_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_22_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_22_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_23_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_23_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_24_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_24_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_25_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_25_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_26_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_26_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_27_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_27_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_28_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_28_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_29_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_29_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_30_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_30_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_31_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_in_31_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_0_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_0_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_1_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_1_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_2_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_2_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_3_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_3_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_4_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_4_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_5_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_5_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_6_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_6_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_7_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_7_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_8_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_8_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_9_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_9_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_10_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_10_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_11_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_11_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_12_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_12_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_13_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_13_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_14_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_14_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_15_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_15_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_16_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_16_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_17_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_17_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_18_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_18_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_19_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_19_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_20_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_20_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_21_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_21_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_22_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_22_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_23_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_23_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_24_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_24_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_25_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_25_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_26_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_26_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_27_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_27_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_28_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_28_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_29_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_29_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_30_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_30_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_31_Re; // @[FFTDesigns.scala 3442:28]
  wire [31:0] FFT_sr_v2_nrv_34_io_out_31_Im; // @[FFTDesigns.scala 3442:28]
  wire [31:0] PermutationsBasic_io_in_0_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_0_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_1_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_1_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_2_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_2_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_3_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_3_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_4_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_4_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_5_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_5_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_6_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_6_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_7_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_7_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_8_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_8_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_9_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_9_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_10_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_10_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_11_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_11_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_12_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_12_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_13_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_13_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_14_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_14_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_15_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_15_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_16_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_16_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_17_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_17_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_18_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_18_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_19_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_19_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_20_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_20_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_21_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_21_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_22_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_22_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_23_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_23_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_24_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_24_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_25_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_25_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_26_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_26_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_27_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_27_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_28_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_28_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_29_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_29_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_30_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_30_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_31_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_31_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_32_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_32_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_33_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_33_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_34_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_34_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_35_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_35_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_36_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_36_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_37_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_37_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_38_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_38_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_39_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_39_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_40_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_40_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_41_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_41_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_42_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_42_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_43_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_43_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_44_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_44_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_45_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_45_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_46_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_46_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_47_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_47_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_48_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_48_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_49_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_49_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_50_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_50_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_51_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_51_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_52_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_52_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_53_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_53_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_54_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_54_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_55_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_55_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_56_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_56_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_57_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_57_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_58_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_58_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_59_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_59_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_60_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_60_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_61_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_61_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_62_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_62_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_63_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_63_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_64_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_64_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_65_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_65_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_66_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_66_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_67_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_67_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_68_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_68_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_69_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_69_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_70_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_70_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_71_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_71_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_72_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_72_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_73_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_73_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_74_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_74_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_75_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_75_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_76_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_76_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_77_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_77_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_78_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_78_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_79_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_79_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_80_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_80_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_81_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_81_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_82_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_82_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_83_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_83_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_84_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_84_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_85_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_85_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_86_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_86_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_87_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_87_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_88_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_88_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_89_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_89_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_90_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_90_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_91_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_91_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_92_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_92_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_93_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_93_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_94_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_94_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_95_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_in_95_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_0_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_0_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_1_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_1_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_2_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_2_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_3_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_3_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_4_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_4_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_5_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_5_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_6_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_6_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_7_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_7_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_8_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_8_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_9_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_9_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_10_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_10_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_11_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_11_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_12_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_12_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_13_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_13_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_14_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_14_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_15_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_15_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_16_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_16_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_17_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_17_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_18_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_18_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_19_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_19_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_20_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_20_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_21_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_21_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_22_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_22_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_23_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_23_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_24_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_24_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_25_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_25_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_26_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_26_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_27_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_27_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_28_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_28_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_29_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_29_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_30_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_30_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_31_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_31_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_32_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_32_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_33_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_33_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_34_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_34_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_35_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_35_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_36_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_36_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_37_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_37_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_38_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_38_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_39_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_39_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_40_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_40_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_41_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_41_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_42_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_42_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_43_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_43_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_44_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_44_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_45_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_45_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_46_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_46_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_47_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_47_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_48_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_48_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_49_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_49_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_50_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_50_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_51_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_51_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_52_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_52_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_53_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_53_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_54_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_54_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_55_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_55_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_56_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_56_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_57_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_57_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_58_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_58_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_59_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_59_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_60_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_60_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_61_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_61_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_62_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_62_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_63_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_63_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_64_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_64_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_65_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_65_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_66_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_66_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_67_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_67_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_68_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_68_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_69_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_69_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_70_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_70_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_71_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_71_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_72_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_72_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_73_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_73_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_74_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_74_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_75_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_75_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_76_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_76_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_77_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_77_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_78_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_78_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_79_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_79_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_80_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_80_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_81_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_81_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_82_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_82_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_83_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_83_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_84_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_84_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_85_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_85_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_86_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_86_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_87_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_87_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_88_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_88_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_89_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_89_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_90_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_90_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_91_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_91_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_92_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_92_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_93_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_93_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_94_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_94_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_95_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_io_out_95_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_1_io_in_0_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_0_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_1_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_1_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_2_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_2_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_3_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_3_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_4_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_4_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_5_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_5_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_6_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_6_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_7_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_7_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_8_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_8_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_9_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_9_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_10_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_10_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_11_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_11_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_12_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_12_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_13_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_13_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_14_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_14_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_15_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_15_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_16_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_16_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_17_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_17_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_18_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_18_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_19_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_19_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_20_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_20_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_21_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_21_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_22_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_22_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_23_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_23_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_24_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_24_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_25_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_25_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_26_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_26_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_27_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_27_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_28_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_28_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_29_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_29_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_30_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_30_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_31_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_31_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_32_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_32_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_33_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_33_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_34_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_34_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_35_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_35_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_36_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_36_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_37_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_37_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_38_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_38_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_39_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_39_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_40_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_40_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_41_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_41_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_42_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_42_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_43_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_43_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_44_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_44_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_45_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_45_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_46_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_46_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_47_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_47_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_48_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_48_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_49_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_49_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_50_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_50_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_51_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_51_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_52_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_52_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_53_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_53_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_54_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_54_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_55_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_55_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_56_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_56_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_57_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_57_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_58_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_58_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_59_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_59_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_60_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_60_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_61_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_61_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_62_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_62_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_63_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_63_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_64_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_64_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_65_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_65_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_66_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_66_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_67_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_67_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_68_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_68_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_69_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_69_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_70_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_70_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_71_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_71_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_72_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_72_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_73_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_73_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_74_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_74_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_75_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_75_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_76_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_76_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_77_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_77_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_78_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_78_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_79_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_79_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_80_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_80_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_81_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_81_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_82_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_82_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_83_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_83_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_84_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_84_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_85_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_85_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_86_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_86_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_87_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_87_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_88_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_88_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_89_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_89_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_90_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_90_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_91_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_91_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_92_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_92_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_93_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_93_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_94_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_94_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_95_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_in_95_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_0_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_0_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_1_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_1_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_2_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_2_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_3_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_3_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_4_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_4_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_5_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_5_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_6_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_6_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_7_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_7_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_8_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_8_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_9_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_9_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_10_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_10_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_11_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_11_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_12_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_12_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_13_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_13_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_14_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_14_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_15_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_15_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_16_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_16_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_17_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_17_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_18_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_18_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_19_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_19_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_20_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_20_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_21_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_21_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_22_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_22_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_23_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_23_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_24_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_24_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_25_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_25_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_26_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_26_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_27_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_27_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_28_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_28_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_29_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_29_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_30_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_30_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_31_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_31_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_32_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_32_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_33_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_33_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_34_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_34_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_35_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_35_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_36_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_36_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_37_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_37_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_38_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_38_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_39_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_39_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_40_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_40_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_41_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_41_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_42_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_42_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_43_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_43_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_44_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_44_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_45_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_45_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_46_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_46_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_47_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_47_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_48_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_48_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_49_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_49_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_50_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_50_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_51_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_51_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_52_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_52_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_53_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_53_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_54_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_54_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_55_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_55_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_56_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_56_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_57_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_57_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_58_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_58_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_59_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_59_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_60_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_60_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_61_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_61_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_62_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_62_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_63_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_63_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_64_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_64_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_65_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_65_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_66_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_66_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_67_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_67_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_68_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_68_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_69_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_69_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_70_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_70_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_71_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_71_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_72_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_72_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_73_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_73_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_74_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_74_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_75_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_75_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_76_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_76_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_77_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_77_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_78_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_78_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_79_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_79_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_80_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_80_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_81_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_81_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_82_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_82_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_83_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_83_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_84_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_84_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_85_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_85_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_86_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_86_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_87_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_87_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_88_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_88_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_89_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_89_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_90_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_90_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_91_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_91_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_92_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_92_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_93_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_93_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_94_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_94_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_95_Re; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_1_io_out_95_Im; // @[FFTDesigns.scala 3447:27]
  wire [31:0] PermutationsBasic_2_io_in_0_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_0_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_1_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_1_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_2_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_2_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_3_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_3_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_4_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_4_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_5_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_5_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_6_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_6_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_7_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_7_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_8_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_8_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_9_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_9_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_10_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_10_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_11_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_11_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_12_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_12_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_13_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_13_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_14_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_14_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_15_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_15_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_16_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_16_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_17_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_17_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_18_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_18_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_19_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_19_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_20_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_20_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_21_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_21_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_22_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_22_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_23_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_23_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_24_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_24_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_25_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_25_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_26_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_26_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_27_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_27_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_28_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_28_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_29_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_29_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_30_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_30_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_31_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_31_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_32_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_32_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_33_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_33_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_34_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_34_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_35_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_35_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_36_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_36_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_37_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_37_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_38_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_38_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_39_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_39_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_40_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_40_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_41_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_41_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_42_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_42_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_43_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_43_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_44_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_44_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_45_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_45_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_46_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_46_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_47_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_47_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_48_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_48_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_49_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_49_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_50_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_50_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_51_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_51_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_52_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_52_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_53_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_53_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_54_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_54_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_55_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_55_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_56_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_56_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_57_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_57_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_58_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_58_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_59_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_59_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_60_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_60_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_61_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_61_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_62_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_62_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_63_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_63_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_64_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_64_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_65_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_65_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_66_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_66_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_67_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_67_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_68_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_68_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_69_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_69_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_70_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_70_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_71_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_71_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_72_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_72_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_73_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_73_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_74_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_74_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_75_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_75_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_76_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_76_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_77_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_77_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_78_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_78_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_79_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_79_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_80_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_80_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_81_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_81_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_82_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_82_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_83_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_83_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_84_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_84_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_85_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_85_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_86_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_86_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_87_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_87_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_88_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_88_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_89_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_89_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_90_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_90_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_91_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_91_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_92_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_92_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_93_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_93_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_94_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_94_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_95_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_in_95_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_0_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_0_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_1_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_1_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_2_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_2_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_3_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_3_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_4_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_4_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_5_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_5_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_6_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_6_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_7_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_7_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_8_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_8_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_9_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_9_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_10_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_10_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_11_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_11_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_12_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_12_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_13_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_13_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_14_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_14_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_15_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_15_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_16_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_16_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_17_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_17_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_18_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_18_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_19_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_19_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_20_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_20_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_21_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_21_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_22_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_22_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_23_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_23_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_24_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_24_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_25_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_25_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_26_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_26_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_27_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_27_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_28_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_28_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_29_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_29_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_30_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_30_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_31_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_31_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_32_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_32_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_33_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_33_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_34_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_34_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_35_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_35_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_36_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_36_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_37_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_37_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_38_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_38_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_39_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_39_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_40_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_40_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_41_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_41_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_42_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_42_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_43_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_43_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_44_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_44_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_45_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_45_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_46_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_46_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_47_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_47_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_48_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_48_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_49_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_49_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_50_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_50_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_51_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_51_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_52_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_52_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_53_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_53_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_54_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_54_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_55_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_55_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_56_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_56_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_57_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_57_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_58_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_58_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_59_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_59_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_60_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_60_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_61_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_61_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_62_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_62_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_63_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_63_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_64_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_64_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_65_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_65_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_66_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_66_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_67_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_67_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_68_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_68_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_69_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_69_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_70_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_70_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_71_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_71_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_72_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_72_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_73_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_73_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_74_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_74_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_75_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_75_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_76_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_76_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_77_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_77_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_78_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_78_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_79_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_79_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_80_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_80_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_81_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_81_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_82_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_82_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_83_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_83_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_84_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_84_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_85_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_85_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_86_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_86_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_87_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_87_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_88_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_88_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_89_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_89_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_90_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_90_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_91_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_91_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_92_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_92_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_93_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_93_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_94_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_94_Im; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_95_Re; // @[FFTDesigns.scala 3450:27]
  wire [31:0] PermutationsBasic_2_io_out_95_Im; // @[FFTDesigns.scala 3450:27]
  wire  TwiddleFactors_mr_clock; // @[FFTDesigns.scala 3454:29]
  wire  TwiddleFactors_mr_reset; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_0_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_0_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_1_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_1_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_2_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_2_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_3_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_3_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_4_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_4_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_5_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_5_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_6_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_6_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_7_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_7_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_8_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_8_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_9_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_9_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_10_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_10_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_11_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_11_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_12_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_12_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_13_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_13_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_14_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_14_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_15_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_15_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_16_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_16_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_17_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_17_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_18_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_18_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_19_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_19_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_20_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_20_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_21_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_21_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_22_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_22_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_23_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_23_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_24_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_24_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_25_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_25_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_26_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_26_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_27_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_27_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_28_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_28_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_29_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_29_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_30_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_30_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_31_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_31_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_32_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_32_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_33_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_33_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_34_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_34_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_35_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_35_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_36_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_36_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_37_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_37_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_38_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_38_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_39_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_39_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_40_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_40_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_41_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_41_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_42_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_42_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_43_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_43_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_44_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_44_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_45_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_45_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_46_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_46_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_47_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_47_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_48_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_48_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_49_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_49_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_50_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_50_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_51_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_51_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_52_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_52_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_53_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_53_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_54_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_54_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_55_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_55_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_56_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_56_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_57_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_57_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_58_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_58_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_59_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_59_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_60_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_60_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_61_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_61_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_62_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_62_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_63_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_63_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_64_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_64_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_65_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_65_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_66_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_66_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_67_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_67_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_68_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_68_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_69_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_69_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_70_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_70_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_71_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_71_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_72_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_72_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_73_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_73_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_74_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_74_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_75_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_75_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_76_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_76_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_77_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_77_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_78_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_78_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_79_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_79_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_80_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_80_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_81_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_81_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_82_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_82_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_83_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_83_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_84_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_84_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_85_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_85_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_86_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_86_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_87_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_87_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_88_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_88_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_89_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_89_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_90_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_90_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_91_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_91_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_92_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_92_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_93_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_93_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_94_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_94_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_95_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_in_95_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_0_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_0_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_1_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_1_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_2_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_2_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_3_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_3_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_4_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_4_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_5_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_5_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_6_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_6_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_7_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_7_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_8_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_8_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_9_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_9_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_10_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_10_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_11_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_11_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_12_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_12_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_13_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_13_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_14_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_14_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_15_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_15_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_16_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_16_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_17_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_17_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_18_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_18_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_19_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_19_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_20_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_20_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_21_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_21_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_22_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_22_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_23_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_23_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_24_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_24_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_25_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_25_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_26_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_26_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_27_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_27_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_28_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_28_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_29_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_29_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_30_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_30_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_31_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_31_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_32_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_32_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_33_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_33_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_34_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_34_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_35_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_35_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_36_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_36_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_37_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_37_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_38_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_38_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_39_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_39_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_40_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_40_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_41_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_41_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_42_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_42_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_43_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_43_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_44_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_44_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_45_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_45_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_46_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_46_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_47_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_47_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_48_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_48_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_49_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_49_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_50_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_50_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_51_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_51_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_52_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_52_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_53_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_53_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_54_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_54_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_55_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_55_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_56_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_56_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_57_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_57_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_58_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_58_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_59_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_59_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_60_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_60_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_61_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_61_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_62_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_62_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_63_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_63_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_64_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_64_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_65_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_65_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_66_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_66_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_67_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_67_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_68_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_68_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_69_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_69_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_70_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_70_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_71_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_71_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_72_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_72_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_73_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_73_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_74_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_74_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_75_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_75_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_76_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_76_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_77_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_77_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_78_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_78_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_79_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_79_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_80_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_80_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_81_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_81_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_82_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_82_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_83_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_83_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_84_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_84_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_85_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_85_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_86_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_86_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_87_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_87_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_88_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_88_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_89_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_89_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_90_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_90_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_91_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_91_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_92_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_92_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_93_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_93_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_94_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_94_Im; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_95_Re; // @[FFTDesigns.scala 3454:29]
  wire [31:0] TwiddleFactors_mr_io_out_95_Im; // @[FFTDesigns.scala 3454:29]
  reg  regdelays_0; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_1; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_2; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_3; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_4; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_5; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_6; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_7; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_8; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_9; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_10; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_11; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_12; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_13; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_14; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_15; // @[FFTDesigns.scala 3427:28]
  reg  regdelays_16; // @[FFTDesigns.scala 3427:28]
  reg  out_regdelay; // @[FFTDesigns.scala 3435:31]
  reg [31:0] out_results_0_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_0_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_1_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_1_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_2_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_2_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_3_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_3_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_4_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_4_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_5_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_5_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_6_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_6_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_7_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_7_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_8_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_8_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_9_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_9_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_10_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_10_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_11_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_11_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_12_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_12_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_13_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_13_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_14_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_14_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_15_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_15_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_16_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_16_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_17_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_17_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_18_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_18_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_19_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_19_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_20_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_20_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_21_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_21_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_22_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_22_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_23_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_23_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_24_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_24_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_25_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_25_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_26_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_26_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_27_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_27_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_28_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_28_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_29_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_29_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_30_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_30_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_31_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_31_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_32_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_32_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_33_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_33_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_34_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_34_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_35_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_35_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_36_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_36_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_37_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_37_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_38_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_38_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_39_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_39_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_40_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_40_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_41_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_41_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_42_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_42_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_43_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_43_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_44_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_44_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_45_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_45_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_46_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_46_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_47_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_47_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_48_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_48_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_49_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_49_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_50_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_50_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_51_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_51_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_52_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_52_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_53_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_53_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_54_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_54_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_55_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_55_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_56_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_56_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_57_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_57_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_58_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_58_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_59_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_59_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_60_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_60_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_61_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_61_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_62_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_62_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_63_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_63_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_64_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_64_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_65_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_65_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_66_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_66_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_67_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_67_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_68_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_68_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_69_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_69_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_70_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_70_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_71_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_71_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_72_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_72_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_73_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_73_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_74_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_74_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_75_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_75_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_76_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_76_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_77_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_77_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_78_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_78_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_79_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_79_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_80_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_80_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_81_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_81_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_82_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_82_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_83_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_83_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_84_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_84_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_85_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_85_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_86_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_86_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_87_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_87_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_88_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_88_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_89_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_89_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_90_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_90_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_91_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_91_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_92_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_92_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_93_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_93_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_94_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_94_Im; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_95_Re; // @[FFTDesigns.scala 3463:30]
  reg [31:0] out_results_95_Im; // @[FFTDesigns.scala 3463:30]
  FFT_sr_v2_nrv FFT_sr_v2_nrv ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_clock),
    .reset(FFT_sr_v2_nrv_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_1 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_1_clock),
    .reset(FFT_sr_v2_nrv_1_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_1_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_1_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_1_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_1_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_1_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_1_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_1_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_1_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_1_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_1_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_1_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_1_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_2 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_2_clock),
    .reset(FFT_sr_v2_nrv_2_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_2_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_2_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_2_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_2_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_2_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_2_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_2_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_2_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_2_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_2_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_2_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_2_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_3 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_3_clock),
    .reset(FFT_sr_v2_nrv_3_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_3_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_3_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_3_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_3_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_3_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_3_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_3_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_3_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_3_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_3_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_3_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_3_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_4 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_4_clock),
    .reset(FFT_sr_v2_nrv_4_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_4_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_4_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_4_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_4_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_4_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_4_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_4_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_4_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_4_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_4_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_4_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_4_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_5 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_5_clock),
    .reset(FFT_sr_v2_nrv_5_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_5_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_5_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_5_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_5_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_5_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_5_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_5_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_5_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_5_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_5_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_5_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_5_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_6 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_6_clock),
    .reset(FFT_sr_v2_nrv_6_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_6_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_6_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_6_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_6_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_6_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_6_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_6_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_6_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_6_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_6_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_6_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_6_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_7 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_7_clock),
    .reset(FFT_sr_v2_nrv_7_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_7_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_7_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_7_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_7_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_7_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_7_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_7_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_7_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_7_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_7_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_7_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_7_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_8 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_8_clock),
    .reset(FFT_sr_v2_nrv_8_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_8_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_8_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_8_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_8_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_8_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_8_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_8_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_8_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_8_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_8_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_8_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_8_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_9 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_9_clock),
    .reset(FFT_sr_v2_nrv_9_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_9_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_9_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_9_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_9_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_9_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_9_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_9_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_9_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_9_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_9_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_9_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_9_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_10 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_10_clock),
    .reset(FFT_sr_v2_nrv_10_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_10_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_10_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_10_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_10_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_10_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_10_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_10_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_10_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_10_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_10_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_10_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_10_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_11 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_11_clock),
    .reset(FFT_sr_v2_nrv_11_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_11_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_11_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_11_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_11_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_11_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_11_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_11_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_11_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_11_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_11_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_11_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_11_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_12 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_12_clock),
    .reset(FFT_sr_v2_nrv_12_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_12_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_12_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_12_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_12_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_12_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_12_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_12_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_12_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_12_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_12_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_12_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_12_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_13 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_13_clock),
    .reset(FFT_sr_v2_nrv_13_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_13_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_13_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_13_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_13_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_13_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_13_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_13_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_13_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_13_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_13_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_13_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_13_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_14 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_14_clock),
    .reset(FFT_sr_v2_nrv_14_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_14_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_14_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_14_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_14_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_14_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_14_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_14_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_14_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_14_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_14_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_14_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_14_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_15 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_15_clock),
    .reset(FFT_sr_v2_nrv_15_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_15_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_15_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_15_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_15_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_15_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_15_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_15_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_15_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_15_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_15_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_15_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_15_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_16 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_16_clock),
    .reset(FFT_sr_v2_nrv_16_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_16_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_16_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_16_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_16_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_16_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_16_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_16_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_16_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_16_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_16_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_16_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_16_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_17 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_17_clock),
    .reset(FFT_sr_v2_nrv_17_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_17_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_17_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_17_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_17_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_17_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_17_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_17_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_17_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_17_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_17_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_17_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_17_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_18 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_18_clock),
    .reset(FFT_sr_v2_nrv_18_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_18_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_18_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_18_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_18_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_18_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_18_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_18_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_18_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_18_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_18_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_18_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_18_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_19 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_19_clock),
    .reset(FFT_sr_v2_nrv_19_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_19_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_19_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_19_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_19_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_19_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_19_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_19_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_19_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_19_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_19_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_19_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_19_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_20 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_20_clock),
    .reset(FFT_sr_v2_nrv_20_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_20_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_20_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_20_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_20_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_20_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_20_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_20_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_20_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_20_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_20_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_20_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_20_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_21 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_21_clock),
    .reset(FFT_sr_v2_nrv_21_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_21_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_21_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_21_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_21_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_21_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_21_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_21_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_21_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_21_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_21_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_21_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_21_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_22 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_22_clock),
    .reset(FFT_sr_v2_nrv_22_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_22_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_22_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_22_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_22_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_22_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_22_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_22_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_22_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_22_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_22_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_22_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_22_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_23 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_23_clock),
    .reset(FFT_sr_v2_nrv_23_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_23_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_23_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_23_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_23_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_23_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_23_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_23_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_23_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_23_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_23_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_23_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_23_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_24 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_24_clock),
    .reset(FFT_sr_v2_nrv_24_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_24_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_24_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_24_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_24_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_24_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_24_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_24_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_24_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_24_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_24_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_24_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_24_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_25 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_25_clock),
    .reset(FFT_sr_v2_nrv_25_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_25_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_25_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_25_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_25_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_25_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_25_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_25_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_25_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_25_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_25_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_25_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_25_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_26 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_26_clock),
    .reset(FFT_sr_v2_nrv_26_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_26_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_26_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_26_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_26_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_26_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_26_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_26_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_26_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_26_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_26_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_26_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_26_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_27 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_27_clock),
    .reset(FFT_sr_v2_nrv_27_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_27_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_27_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_27_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_27_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_27_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_27_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_27_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_27_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_27_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_27_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_27_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_27_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_28 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_28_clock),
    .reset(FFT_sr_v2_nrv_28_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_28_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_28_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_28_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_28_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_28_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_28_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_28_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_28_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_28_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_28_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_28_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_28_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_29 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_29_clock),
    .reset(FFT_sr_v2_nrv_29_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_29_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_29_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_29_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_29_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_29_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_29_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_29_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_29_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_29_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_29_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_29_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_29_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_30 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_30_clock),
    .reset(FFT_sr_v2_nrv_30_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_30_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_30_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_30_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_30_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_30_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_30_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_30_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_30_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_30_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_30_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_30_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_30_io_out_2_Im)
  );
  FFT_sr_v2_nrv FFT_sr_v2_nrv_31 ( // @[FFTDesigns.scala 3438:28]
    .clock(FFT_sr_v2_nrv_31_clock),
    .reset(FFT_sr_v2_nrv_31_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_31_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_31_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_31_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_31_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_31_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_31_io_in_2_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_31_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_31_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_31_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_31_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_31_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_31_io_out_2_Im)
  );
  FFT_sr_v2_nrv_32 FFT_sr_v2_nrv_32 ( // @[FFTDesigns.scala 3442:28]
    .clock(FFT_sr_v2_nrv_32_clock),
    .reset(FFT_sr_v2_nrv_32_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_32_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_32_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_32_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_32_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_32_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_32_io_in_2_Im),
    .io_in_3_Re(FFT_sr_v2_nrv_32_io_in_3_Re),
    .io_in_3_Im(FFT_sr_v2_nrv_32_io_in_3_Im),
    .io_in_4_Re(FFT_sr_v2_nrv_32_io_in_4_Re),
    .io_in_4_Im(FFT_sr_v2_nrv_32_io_in_4_Im),
    .io_in_5_Re(FFT_sr_v2_nrv_32_io_in_5_Re),
    .io_in_5_Im(FFT_sr_v2_nrv_32_io_in_5_Im),
    .io_in_6_Re(FFT_sr_v2_nrv_32_io_in_6_Re),
    .io_in_6_Im(FFT_sr_v2_nrv_32_io_in_6_Im),
    .io_in_7_Re(FFT_sr_v2_nrv_32_io_in_7_Re),
    .io_in_7_Im(FFT_sr_v2_nrv_32_io_in_7_Im),
    .io_in_8_Re(FFT_sr_v2_nrv_32_io_in_8_Re),
    .io_in_8_Im(FFT_sr_v2_nrv_32_io_in_8_Im),
    .io_in_9_Re(FFT_sr_v2_nrv_32_io_in_9_Re),
    .io_in_9_Im(FFT_sr_v2_nrv_32_io_in_9_Im),
    .io_in_10_Re(FFT_sr_v2_nrv_32_io_in_10_Re),
    .io_in_10_Im(FFT_sr_v2_nrv_32_io_in_10_Im),
    .io_in_11_Re(FFT_sr_v2_nrv_32_io_in_11_Re),
    .io_in_11_Im(FFT_sr_v2_nrv_32_io_in_11_Im),
    .io_in_12_Re(FFT_sr_v2_nrv_32_io_in_12_Re),
    .io_in_12_Im(FFT_sr_v2_nrv_32_io_in_12_Im),
    .io_in_13_Re(FFT_sr_v2_nrv_32_io_in_13_Re),
    .io_in_13_Im(FFT_sr_v2_nrv_32_io_in_13_Im),
    .io_in_14_Re(FFT_sr_v2_nrv_32_io_in_14_Re),
    .io_in_14_Im(FFT_sr_v2_nrv_32_io_in_14_Im),
    .io_in_15_Re(FFT_sr_v2_nrv_32_io_in_15_Re),
    .io_in_15_Im(FFT_sr_v2_nrv_32_io_in_15_Im),
    .io_in_16_Re(FFT_sr_v2_nrv_32_io_in_16_Re),
    .io_in_16_Im(FFT_sr_v2_nrv_32_io_in_16_Im),
    .io_in_17_Re(FFT_sr_v2_nrv_32_io_in_17_Re),
    .io_in_17_Im(FFT_sr_v2_nrv_32_io_in_17_Im),
    .io_in_18_Re(FFT_sr_v2_nrv_32_io_in_18_Re),
    .io_in_18_Im(FFT_sr_v2_nrv_32_io_in_18_Im),
    .io_in_19_Re(FFT_sr_v2_nrv_32_io_in_19_Re),
    .io_in_19_Im(FFT_sr_v2_nrv_32_io_in_19_Im),
    .io_in_20_Re(FFT_sr_v2_nrv_32_io_in_20_Re),
    .io_in_20_Im(FFT_sr_v2_nrv_32_io_in_20_Im),
    .io_in_21_Re(FFT_sr_v2_nrv_32_io_in_21_Re),
    .io_in_21_Im(FFT_sr_v2_nrv_32_io_in_21_Im),
    .io_in_22_Re(FFT_sr_v2_nrv_32_io_in_22_Re),
    .io_in_22_Im(FFT_sr_v2_nrv_32_io_in_22_Im),
    .io_in_23_Re(FFT_sr_v2_nrv_32_io_in_23_Re),
    .io_in_23_Im(FFT_sr_v2_nrv_32_io_in_23_Im),
    .io_in_24_Re(FFT_sr_v2_nrv_32_io_in_24_Re),
    .io_in_24_Im(FFT_sr_v2_nrv_32_io_in_24_Im),
    .io_in_25_Re(FFT_sr_v2_nrv_32_io_in_25_Re),
    .io_in_25_Im(FFT_sr_v2_nrv_32_io_in_25_Im),
    .io_in_26_Re(FFT_sr_v2_nrv_32_io_in_26_Re),
    .io_in_26_Im(FFT_sr_v2_nrv_32_io_in_26_Im),
    .io_in_27_Re(FFT_sr_v2_nrv_32_io_in_27_Re),
    .io_in_27_Im(FFT_sr_v2_nrv_32_io_in_27_Im),
    .io_in_28_Re(FFT_sr_v2_nrv_32_io_in_28_Re),
    .io_in_28_Im(FFT_sr_v2_nrv_32_io_in_28_Im),
    .io_in_29_Re(FFT_sr_v2_nrv_32_io_in_29_Re),
    .io_in_29_Im(FFT_sr_v2_nrv_32_io_in_29_Im),
    .io_in_30_Re(FFT_sr_v2_nrv_32_io_in_30_Re),
    .io_in_30_Im(FFT_sr_v2_nrv_32_io_in_30_Im),
    .io_in_31_Re(FFT_sr_v2_nrv_32_io_in_31_Re),
    .io_in_31_Im(FFT_sr_v2_nrv_32_io_in_31_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_32_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_32_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_32_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_32_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_32_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_32_io_out_2_Im),
    .io_out_3_Re(FFT_sr_v2_nrv_32_io_out_3_Re),
    .io_out_3_Im(FFT_sr_v2_nrv_32_io_out_3_Im),
    .io_out_4_Re(FFT_sr_v2_nrv_32_io_out_4_Re),
    .io_out_4_Im(FFT_sr_v2_nrv_32_io_out_4_Im),
    .io_out_5_Re(FFT_sr_v2_nrv_32_io_out_5_Re),
    .io_out_5_Im(FFT_sr_v2_nrv_32_io_out_5_Im),
    .io_out_6_Re(FFT_sr_v2_nrv_32_io_out_6_Re),
    .io_out_6_Im(FFT_sr_v2_nrv_32_io_out_6_Im),
    .io_out_7_Re(FFT_sr_v2_nrv_32_io_out_7_Re),
    .io_out_7_Im(FFT_sr_v2_nrv_32_io_out_7_Im),
    .io_out_8_Re(FFT_sr_v2_nrv_32_io_out_8_Re),
    .io_out_8_Im(FFT_sr_v2_nrv_32_io_out_8_Im),
    .io_out_9_Re(FFT_sr_v2_nrv_32_io_out_9_Re),
    .io_out_9_Im(FFT_sr_v2_nrv_32_io_out_9_Im),
    .io_out_10_Re(FFT_sr_v2_nrv_32_io_out_10_Re),
    .io_out_10_Im(FFT_sr_v2_nrv_32_io_out_10_Im),
    .io_out_11_Re(FFT_sr_v2_nrv_32_io_out_11_Re),
    .io_out_11_Im(FFT_sr_v2_nrv_32_io_out_11_Im),
    .io_out_12_Re(FFT_sr_v2_nrv_32_io_out_12_Re),
    .io_out_12_Im(FFT_sr_v2_nrv_32_io_out_12_Im),
    .io_out_13_Re(FFT_sr_v2_nrv_32_io_out_13_Re),
    .io_out_13_Im(FFT_sr_v2_nrv_32_io_out_13_Im),
    .io_out_14_Re(FFT_sr_v2_nrv_32_io_out_14_Re),
    .io_out_14_Im(FFT_sr_v2_nrv_32_io_out_14_Im),
    .io_out_15_Re(FFT_sr_v2_nrv_32_io_out_15_Re),
    .io_out_15_Im(FFT_sr_v2_nrv_32_io_out_15_Im),
    .io_out_16_Re(FFT_sr_v2_nrv_32_io_out_16_Re),
    .io_out_16_Im(FFT_sr_v2_nrv_32_io_out_16_Im),
    .io_out_17_Re(FFT_sr_v2_nrv_32_io_out_17_Re),
    .io_out_17_Im(FFT_sr_v2_nrv_32_io_out_17_Im),
    .io_out_18_Re(FFT_sr_v2_nrv_32_io_out_18_Re),
    .io_out_18_Im(FFT_sr_v2_nrv_32_io_out_18_Im),
    .io_out_19_Re(FFT_sr_v2_nrv_32_io_out_19_Re),
    .io_out_19_Im(FFT_sr_v2_nrv_32_io_out_19_Im),
    .io_out_20_Re(FFT_sr_v2_nrv_32_io_out_20_Re),
    .io_out_20_Im(FFT_sr_v2_nrv_32_io_out_20_Im),
    .io_out_21_Re(FFT_sr_v2_nrv_32_io_out_21_Re),
    .io_out_21_Im(FFT_sr_v2_nrv_32_io_out_21_Im),
    .io_out_22_Re(FFT_sr_v2_nrv_32_io_out_22_Re),
    .io_out_22_Im(FFT_sr_v2_nrv_32_io_out_22_Im),
    .io_out_23_Re(FFT_sr_v2_nrv_32_io_out_23_Re),
    .io_out_23_Im(FFT_sr_v2_nrv_32_io_out_23_Im),
    .io_out_24_Re(FFT_sr_v2_nrv_32_io_out_24_Re),
    .io_out_24_Im(FFT_sr_v2_nrv_32_io_out_24_Im),
    .io_out_25_Re(FFT_sr_v2_nrv_32_io_out_25_Re),
    .io_out_25_Im(FFT_sr_v2_nrv_32_io_out_25_Im),
    .io_out_26_Re(FFT_sr_v2_nrv_32_io_out_26_Re),
    .io_out_26_Im(FFT_sr_v2_nrv_32_io_out_26_Im),
    .io_out_27_Re(FFT_sr_v2_nrv_32_io_out_27_Re),
    .io_out_27_Im(FFT_sr_v2_nrv_32_io_out_27_Im),
    .io_out_28_Re(FFT_sr_v2_nrv_32_io_out_28_Re),
    .io_out_28_Im(FFT_sr_v2_nrv_32_io_out_28_Im),
    .io_out_29_Re(FFT_sr_v2_nrv_32_io_out_29_Re),
    .io_out_29_Im(FFT_sr_v2_nrv_32_io_out_29_Im),
    .io_out_30_Re(FFT_sr_v2_nrv_32_io_out_30_Re),
    .io_out_30_Im(FFT_sr_v2_nrv_32_io_out_30_Im),
    .io_out_31_Re(FFT_sr_v2_nrv_32_io_out_31_Re),
    .io_out_31_Im(FFT_sr_v2_nrv_32_io_out_31_Im)
  );
  FFT_sr_v2_nrv_32 FFT_sr_v2_nrv_33 ( // @[FFTDesigns.scala 3442:28]
    .clock(FFT_sr_v2_nrv_33_clock),
    .reset(FFT_sr_v2_nrv_33_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_33_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_33_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_33_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_33_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_33_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_33_io_in_2_Im),
    .io_in_3_Re(FFT_sr_v2_nrv_33_io_in_3_Re),
    .io_in_3_Im(FFT_sr_v2_nrv_33_io_in_3_Im),
    .io_in_4_Re(FFT_sr_v2_nrv_33_io_in_4_Re),
    .io_in_4_Im(FFT_sr_v2_nrv_33_io_in_4_Im),
    .io_in_5_Re(FFT_sr_v2_nrv_33_io_in_5_Re),
    .io_in_5_Im(FFT_sr_v2_nrv_33_io_in_5_Im),
    .io_in_6_Re(FFT_sr_v2_nrv_33_io_in_6_Re),
    .io_in_6_Im(FFT_sr_v2_nrv_33_io_in_6_Im),
    .io_in_7_Re(FFT_sr_v2_nrv_33_io_in_7_Re),
    .io_in_7_Im(FFT_sr_v2_nrv_33_io_in_7_Im),
    .io_in_8_Re(FFT_sr_v2_nrv_33_io_in_8_Re),
    .io_in_8_Im(FFT_sr_v2_nrv_33_io_in_8_Im),
    .io_in_9_Re(FFT_sr_v2_nrv_33_io_in_9_Re),
    .io_in_9_Im(FFT_sr_v2_nrv_33_io_in_9_Im),
    .io_in_10_Re(FFT_sr_v2_nrv_33_io_in_10_Re),
    .io_in_10_Im(FFT_sr_v2_nrv_33_io_in_10_Im),
    .io_in_11_Re(FFT_sr_v2_nrv_33_io_in_11_Re),
    .io_in_11_Im(FFT_sr_v2_nrv_33_io_in_11_Im),
    .io_in_12_Re(FFT_sr_v2_nrv_33_io_in_12_Re),
    .io_in_12_Im(FFT_sr_v2_nrv_33_io_in_12_Im),
    .io_in_13_Re(FFT_sr_v2_nrv_33_io_in_13_Re),
    .io_in_13_Im(FFT_sr_v2_nrv_33_io_in_13_Im),
    .io_in_14_Re(FFT_sr_v2_nrv_33_io_in_14_Re),
    .io_in_14_Im(FFT_sr_v2_nrv_33_io_in_14_Im),
    .io_in_15_Re(FFT_sr_v2_nrv_33_io_in_15_Re),
    .io_in_15_Im(FFT_sr_v2_nrv_33_io_in_15_Im),
    .io_in_16_Re(FFT_sr_v2_nrv_33_io_in_16_Re),
    .io_in_16_Im(FFT_sr_v2_nrv_33_io_in_16_Im),
    .io_in_17_Re(FFT_sr_v2_nrv_33_io_in_17_Re),
    .io_in_17_Im(FFT_sr_v2_nrv_33_io_in_17_Im),
    .io_in_18_Re(FFT_sr_v2_nrv_33_io_in_18_Re),
    .io_in_18_Im(FFT_sr_v2_nrv_33_io_in_18_Im),
    .io_in_19_Re(FFT_sr_v2_nrv_33_io_in_19_Re),
    .io_in_19_Im(FFT_sr_v2_nrv_33_io_in_19_Im),
    .io_in_20_Re(FFT_sr_v2_nrv_33_io_in_20_Re),
    .io_in_20_Im(FFT_sr_v2_nrv_33_io_in_20_Im),
    .io_in_21_Re(FFT_sr_v2_nrv_33_io_in_21_Re),
    .io_in_21_Im(FFT_sr_v2_nrv_33_io_in_21_Im),
    .io_in_22_Re(FFT_sr_v2_nrv_33_io_in_22_Re),
    .io_in_22_Im(FFT_sr_v2_nrv_33_io_in_22_Im),
    .io_in_23_Re(FFT_sr_v2_nrv_33_io_in_23_Re),
    .io_in_23_Im(FFT_sr_v2_nrv_33_io_in_23_Im),
    .io_in_24_Re(FFT_sr_v2_nrv_33_io_in_24_Re),
    .io_in_24_Im(FFT_sr_v2_nrv_33_io_in_24_Im),
    .io_in_25_Re(FFT_sr_v2_nrv_33_io_in_25_Re),
    .io_in_25_Im(FFT_sr_v2_nrv_33_io_in_25_Im),
    .io_in_26_Re(FFT_sr_v2_nrv_33_io_in_26_Re),
    .io_in_26_Im(FFT_sr_v2_nrv_33_io_in_26_Im),
    .io_in_27_Re(FFT_sr_v2_nrv_33_io_in_27_Re),
    .io_in_27_Im(FFT_sr_v2_nrv_33_io_in_27_Im),
    .io_in_28_Re(FFT_sr_v2_nrv_33_io_in_28_Re),
    .io_in_28_Im(FFT_sr_v2_nrv_33_io_in_28_Im),
    .io_in_29_Re(FFT_sr_v2_nrv_33_io_in_29_Re),
    .io_in_29_Im(FFT_sr_v2_nrv_33_io_in_29_Im),
    .io_in_30_Re(FFT_sr_v2_nrv_33_io_in_30_Re),
    .io_in_30_Im(FFT_sr_v2_nrv_33_io_in_30_Im),
    .io_in_31_Re(FFT_sr_v2_nrv_33_io_in_31_Re),
    .io_in_31_Im(FFT_sr_v2_nrv_33_io_in_31_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_33_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_33_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_33_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_33_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_33_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_33_io_out_2_Im),
    .io_out_3_Re(FFT_sr_v2_nrv_33_io_out_3_Re),
    .io_out_3_Im(FFT_sr_v2_nrv_33_io_out_3_Im),
    .io_out_4_Re(FFT_sr_v2_nrv_33_io_out_4_Re),
    .io_out_4_Im(FFT_sr_v2_nrv_33_io_out_4_Im),
    .io_out_5_Re(FFT_sr_v2_nrv_33_io_out_5_Re),
    .io_out_5_Im(FFT_sr_v2_nrv_33_io_out_5_Im),
    .io_out_6_Re(FFT_sr_v2_nrv_33_io_out_6_Re),
    .io_out_6_Im(FFT_sr_v2_nrv_33_io_out_6_Im),
    .io_out_7_Re(FFT_sr_v2_nrv_33_io_out_7_Re),
    .io_out_7_Im(FFT_sr_v2_nrv_33_io_out_7_Im),
    .io_out_8_Re(FFT_sr_v2_nrv_33_io_out_8_Re),
    .io_out_8_Im(FFT_sr_v2_nrv_33_io_out_8_Im),
    .io_out_9_Re(FFT_sr_v2_nrv_33_io_out_9_Re),
    .io_out_9_Im(FFT_sr_v2_nrv_33_io_out_9_Im),
    .io_out_10_Re(FFT_sr_v2_nrv_33_io_out_10_Re),
    .io_out_10_Im(FFT_sr_v2_nrv_33_io_out_10_Im),
    .io_out_11_Re(FFT_sr_v2_nrv_33_io_out_11_Re),
    .io_out_11_Im(FFT_sr_v2_nrv_33_io_out_11_Im),
    .io_out_12_Re(FFT_sr_v2_nrv_33_io_out_12_Re),
    .io_out_12_Im(FFT_sr_v2_nrv_33_io_out_12_Im),
    .io_out_13_Re(FFT_sr_v2_nrv_33_io_out_13_Re),
    .io_out_13_Im(FFT_sr_v2_nrv_33_io_out_13_Im),
    .io_out_14_Re(FFT_sr_v2_nrv_33_io_out_14_Re),
    .io_out_14_Im(FFT_sr_v2_nrv_33_io_out_14_Im),
    .io_out_15_Re(FFT_sr_v2_nrv_33_io_out_15_Re),
    .io_out_15_Im(FFT_sr_v2_nrv_33_io_out_15_Im),
    .io_out_16_Re(FFT_sr_v2_nrv_33_io_out_16_Re),
    .io_out_16_Im(FFT_sr_v2_nrv_33_io_out_16_Im),
    .io_out_17_Re(FFT_sr_v2_nrv_33_io_out_17_Re),
    .io_out_17_Im(FFT_sr_v2_nrv_33_io_out_17_Im),
    .io_out_18_Re(FFT_sr_v2_nrv_33_io_out_18_Re),
    .io_out_18_Im(FFT_sr_v2_nrv_33_io_out_18_Im),
    .io_out_19_Re(FFT_sr_v2_nrv_33_io_out_19_Re),
    .io_out_19_Im(FFT_sr_v2_nrv_33_io_out_19_Im),
    .io_out_20_Re(FFT_sr_v2_nrv_33_io_out_20_Re),
    .io_out_20_Im(FFT_sr_v2_nrv_33_io_out_20_Im),
    .io_out_21_Re(FFT_sr_v2_nrv_33_io_out_21_Re),
    .io_out_21_Im(FFT_sr_v2_nrv_33_io_out_21_Im),
    .io_out_22_Re(FFT_sr_v2_nrv_33_io_out_22_Re),
    .io_out_22_Im(FFT_sr_v2_nrv_33_io_out_22_Im),
    .io_out_23_Re(FFT_sr_v2_nrv_33_io_out_23_Re),
    .io_out_23_Im(FFT_sr_v2_nrv_33_io_out_23_Im),
    .io_out_24_Re(FFT_sr_v2_nrv_33_io_out_24_Re),
    .io_out_24_Im(FFT_sr_v2_nrv_33_io_out_24_Im),
    .io_out_25_Re(FFT_sr_v2_nrv_33_io_out_25_Re),
    .io_out_25_Im(FFT_sr_v2_nrv_33_io_out_25_Im),
    .io_out_26_Re(FFT_sr_v2_nrv_33_io_out_26_Re),
    .io_out_26_Im(FFT_sr_v2_nrv_33_io_out_26_Im),
    .io_out_27_Re(FFT_sr_v2_nrv_33_io_out_27_Re),
    .io_out_27_Im(FFT_sr_v2_nrv_33_io_out_27_Im),
    .io_out_28_Re(FFT_sr_v2_nrv_33_io_out_28_Re),
    .io_out_28_Im(FFT_sr_v2_nrv_33_io_out_28_Im),
    .io_out_29_Re(FFT_sr_v2_nrv_33_io_out_29_Re),
    .io_out_29_Im(FFT_sr_v2_nrv_33_io_out_29_Im),
    .io_out_30_Re(FFT_sr_v2_nrv_33_io_out_30_Re),
    .io_out_30_Im(FFT_sr_v2_nrv_33_io_out_30_Im),
    .io_out_31_Re(FFT_sr_v2_nrv_33_io_out_31_Re),
    .io_out_31_Im(FFT_sr_v2_nrv_33_io_out_31_Im)
  );
  FFT_sr_v2_nrv_32 FFT_sr_v2_nrv_34 ( // @[FFTDesigns.scala 3442:28]
    .clock(FFT_sr_v2_nrv_34_clock),
    .reset(FFT_sr_v2_nrv_34_reset),
    .io_in_0_Re(FFT_sr_v2_nrv_34_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_nrv_34_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_nrv_34_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_nrv_34_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_nrv_34_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_nrv_34_io_in_2_Im),
    .io_in_3_Re(FFT_sr_v2_nrv_34_io_in_3_Re),
    .io_in_3_Im(FFT_sr_v2_nrv_34_io_in_3_Im),
    .io_in_4_Re(FFT_sr_v2_nrv_34_io_in_4_Re),
    .io_in_4_Im(FFT_sr_v2_nrv_34_io_in_4_Im),
    .io_in_5_Re(FFT_sr_v2_nrv_34_io_in_5_Re),
    .io_in_5_Im(FFT_sr_v2_nrv_34_io_in_5_Im),
    .io_in_6_Re(FFT_sr_v2_nrv_34_io_in_6_Re),
    .io_in_6_Im(FFT_sr_v2_nrv_34_io_in_6_Im),
    .io_in_7_Re(FFT_sr_v2_nrv_34_io_in_7_Re),
    .io_in_7_Im(FFT_sr_v2_nrv_34_io_in_7_Im),
    .io_in_8_Re(FFT_sr_v2_nrv_34_io_in_8_Re),
    .io_in_8_Im(FFT_sr_v2_nrv_34_io_in_8_Im),
    .io_in_9_Re(FFT_sr_v2_nrv_34_io_in_9_Re),
    .io_in_9_Im(FFT_sr_v2_nrv_34_io_in_9_Im),
    .io_in_10_Re(FFT_sr_v2_nrv_34_io_in_10_Re),
    .io_in_10_Im(FFT_sr_v2_nrv_34_io_in_10_Im),
    .io_in_11_Re(FFT_sr_v2_nrv_34_io_in_11_Re),
    .io_in_11_Im(FFT_sr_v2_nrv_34_io_in_11_Im),
    .io_in_12_Re(FFT_sr_v2_nrv_34_io_in_12_Re),
    .io_in_12_Im(FFT_sr_v2_nrv_34_io_in_12_Im),
    .io_in_13_Re(FFT_sr_v2_nrv_34_io_in_13_Re),
    .io_in_13_Im(FFT_sr_v2_nrv_34_io_in_13_Im),
    .io_in_14_Re(FFT_sr_v2_nrv_34_io_in_14_Re),
    .io_in_14_Im(FFT_sr_v2_nrv_34_io_in_14_Im),
    .io_in_15_Re(FFT_sr_v2_nrv_34_io_in_15_Re),
    .io_in_15_Im(FFT_sr_v2_nrv_34_io_in_15_Im),
    .io_in_16_Re(FFT_sr_v2_nrv_34_io_in_16_Re),
    .io_in_16_Im(FFT_sr_v2_nrv_34_io_in_16_Im),
    .io_in_17_Re(FFT_sr_v2_nrv_34_io_in_17_Re),
    .io_in_17_Im(FFT_sr_v2_nrv_34_io_in_17_Im),
    .io_in_18_Re(FFT_sr_v2_nrv_34_io_in_18_Re),
    .io_in_18_Im(FFT_sr_v2_nrv_34_io_in_18_Im),
    .io_in_19_Re(FFT_sr_v2_nrv_34_io_in_19_Re),
    .io_in_19_Im(FFT_sr_v2_nrv_34_io_in_19_Im),
    .io_in_20_Re(FFT_sr_v2_nrv_34_io_in_20_Re),
    .io_in_20_Im(FFT_sr_v2_nrv_34_io_in_20_Im),
    .io_in_21_Re(FFT_sr_v2_nrv_34_io_in_21_Re),
    .io_in_21_Im(FFT_sr_v2_nrv_34_io_in_21_Im),
    .io_in_22_Re(FFT_sr_v2_nrv_34_io_in_22_Re),
    .io_in_22_Im(FFT_sr_v2_nrv_34_io_in_22_Im),
    .io_in_23_Re(FFT_sr_v2_nrv_34_io_in_23_Re),
    .io_in_23_Im(FFT_sr_v2_nrv_34_io_in_23_Im),
    .io_in_24_Re(FFT_sr_v2_nrv_34_io_in_24_Re),
    .io_in_24_Im(FFT_sr_v2_nrv_34_io_in_24_Im),
    .io_in_25_Re(FFT_sr_v2_nrv_34_io_in_25_Re),
    .io_in_25_Im(FFT_sr_v2_nrv_34_io_in_25_Im),
    .io_in_26_Re(FFT_sr_v2_nrv_34_io_in_26_Re),
    .io_in_26_Im(FFT_sr_v2_nrv_34_io_in_26_Im),
    .io_in_27_Re(FFT_sr_v2_nrv_34_io_in_27_Re),
    .io_in_27_Im(FFT_sr_v2_nrv_34_io_in_27_Im),
    .io_in_28_Re(FFT_sr_v2_nrv_34_io_in_28_Re),
    .io_in_28_Im(FFT_sr_v2_nrv_34_io_in_28_Im),
    .io_in_29_Re(FFT_sr_v2_nrv_34_io_in_29_Re),
    .io_in_29_Im(FFT_sr_v2_nrv_34_io_in_29_Im),
    .io_in_30_Re(FFT_sr_v2_nrv_34_io_in_30_Re),
    .io_in_30_Im(FFT_sr_v2_nrv_34_io_in_30_Im),
    .io_in_31_Re(FFT_sr_v2_nrv_34_io_in_31_Re),
    .io_in_31_Im(FFT_sr_v2_nrv_34_io_in_31_Im),
    .io_out_0_Re(FFT_sr_v2_nrv_34_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_nrv_34_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_nrv_34_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_nrv_34_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_nrv_34_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_nrv_34_io_out_2_Im),
    .io_out_3_Re(FFT_sr_v2_nrv_34_io_out_3_Re),
    .io_out_3_Im(FFT_sr_v2_nrv_34_io_out_3_Im),
    .io_out_4_Re(FFT_sr_v2_nrv_34_io_out_4_Re),
    .io_out_4_Im(FFT_sr_v2_nrv_34_io_out_4_Im),
    .io_out_5_Re(FFT_sr_v2_nrv_34_io_out_5_Re),
    .io_out_5_Im(FFT_sr_v2_nrv_34_io_out_5_Im),
    .io_out_6_Re(FFT_sr_v2_nrv_34_io_out_6_Re),
    .io_out_6_Im(FFT_sr_v2_nrv_34_io_out_6_Im),
    .io_out_7_Re(FFT_sr_v2_nrv_34_io_out_7_Re),
    .io_out_7_Im(FFT_sr_v2_nrv_34_io_out_7_Im),
    .io_out_8_Re(FFT_sr_v2_nrv_34_io_out_8_Re),
    .io_out_8_Im(FFT_sr_v2_nrv_34_io_out_8_Im),
    .io_out_9_Re(FFT_sr_v2_nrv_34_io_out_9_Re),
    .io_out_9_Im(FFT_sr_v2_nrv_34_io_out_9_Im),
    .io_out_10_Re(FFT_sr_v2_nrv_34_io_out_10_Re),
    .io_out_10_Im(FFT_sr_v2_nrv_34_io_out_10_Im),
    .io_out_11_Re(FFT_sr_v2_nrv_34_io_out_11_Re),
    .io_out_11_Im(FFT_sr_v2_nrv_34_io_out_11_Im),
    .io_out_12_Re(FFT_sr_v2_nrv_34_io_out_12_Re),
    .io_out_12_Im(FFT_sr_v2_nrv_34_io_out_12_Im),
    .io_out_13_Re(FFT_sr_v2_nrv_34_io_out_13_Re),
    .io_out_13_Im(FFT_sr_v2_nrv_34_io_out_13_Im),
    .io_out_14_Re(FFT_sr_v2_nrv_34_io_out_14_Re),
    .io_out_14_Im(FFT_sr_v2_nrv_34_io_out_14_Im),
    .io_out_15_Re(FFT_sr_v2_nrv_34_io_out_15_Re),
    .io_out_15_Im(FFT_sr_v2_nrv_34_io_out_15_Im),
    .io_out_16_Re(FFT_sr_v2_nrv_34_io_out_16_Re),
    .io_out_16_Im(FFT_sr_v2_nrv_34_io_out_16_Im),
    .io_out_17_Re(FFT_sr_v2_nrv_34_io_out_17_Re),
    .io_out_17_Im(FFT_sr_v2_nrv_34_io_out_17_Im),
    .io_out_18_Re(FFT_sr_v2_nrv_34_io_out_18_Re),
    .io_out_18_Im(FFT_sr_v2_nrv_34_io_out_18_Im),
    .io_out_19_Re(FFT_sr_v2_nrv_34_io_out_19_Re),
    .io_out_19_Im(FFT_sr_v2_nrv_34_io_out_19_Im),
    .io_out_20_Re(FFT_sr_v2_nrv_34_io_out_20_Re),
    .io_out_20_Im(FFT_sr_v2_nrv_34_io_out_20_Im),
    .io_out_21_Re(FFT_sr_v2_nrv_34_io_out_21_Re),
    .io_out_21_Im(FFT_sr_v2_nrv_34_io_out_21_Im),
    .io_out_22_Re(FFT_sr_v2_nrv_34_io_out_22_Re),
    .io_out_22_Im(FFT_sr_v2_nrv_34_io_out_22_Im),
    .io_out_23_Re(FFT_sr_v2_nrv_34_io_out_23_Re),
    .io_out_23_Im(FFT_sr_v2_nrv_34_io_out_23_Im),
    .io_out_24_Re(FFT_sr_v2_nrv_34_io_out_24_Re),
    .io_out_24_Im(FFT_sr_v2_nrv_34_io_out_24_Im),
    .io_out_25_Re(FFT_sr_v2_nrv_34_io_out_25_Re),
    .io_out_25_Im(FFT_sr_v2_nrv_34_io_out_25_Im),
    .io_out_26_Re(FFT_sr_v2_nrv_34_io_out_26_Re),
    .io_out_26_Im(FFT_sr_v2_nrv_34_io_out_26_Im),
    .io_out_27_Re(FFT_sr_v2_nrv_34_io_out_27_Re),
    .io_out_27_Im(FFT_sr_v2_nrv_34_io_out_27_Im),
    .io_out_28_Re(FFT_sr_v2_nrv_34_io_out_28_Re),
    .io_out_28_Im(FFT_sr_v2_nrv_34_io_out_28_Im),
    .io_out_29_Re(FFT_sr_v2_nrv_34_io_out_29_Re),
    .io_out_29_Im(FFT_sr_v2_nrv_34_io_out_29_Im),
    .io_out_30_Re(FFT_sr_v2_nrv_34_io_out_30_Re),
    .io_out_30_Im(FFT_sr_v2_nrv_34_io_out_30_Im),
    .io_out_31_Re(FFT_sr_v2_nrv_34_io_out_31_Re),
    .io_out_31_Im(FFT_sr_v2_nrv_34_io_out_31_Im)
  );
  PermutationsBasic_82 PermutationsBasic ( // @[FFTDesigns.scala 3450:27]
    .io_in_0_Re(PermutationsBasic_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_io_in_31_Im),
    .io_in_32_Re(PermutationsBasic_io_in_32_Re),
    .io_in_32_Im(PermutationsBasic_io_in_32_Im),
    .io_in_33_Re(PermutationsBasic_io_in_33_Re),
    .io_in_33_Im(PermutationsBasic_io_in_33_Im),
    .io_in_34_Re(PermutationsBasic_io_in_34_Re),
    .io_in_34_Im(PermutationsBasic_io_in_34_Im),
    .io_in_35_Re(PermutationsBasic_io_in_35_Re),
    .io_in_35_Im(PermutationsBasic_io_in_35_Im),
    .io_in_36_Re(PermutationsBasic_io_in_36_Re),
    .io_in_36_Im(PermutationsBasic_io_in_36_Im),
    .io_in_37_Re(PermutationsBasic_io_in_37_Re),
    .io_in_37_Im(PermutationsBasic_io_in_37_Im),
    .io_in_38_Re(PermutationsBasic_io_in_38_Re),
    .io_in_38_Im(PermutationsBasic_io_in_38_Im),
    .io_in_39_Re(PermutationsBasic_io_in_39_Re),
    .io_in_39_Im(PermutationsBasic_io_in_39_Im),
    .io_in_40_Re(PermutationsBasic_io_in_40_Re),
    .io_in_40_Im(PermutationsBasic_io_in_40_Im),
    .io_in_41_Re(PermutationsBasic_io_in_41_Re),
    .io_in_41_Im(PermutationsBasic_io_in_41_Im),
    .io_in_42_Re(PermutationsBasic_io_in_42_Re),
    .io_in_42_Im(PermutationsBasic_io_in_42_Im),
    .io_in_43_Re(PermutationsBasic_io_in_43_Re),
    .io_in_43_Im(PermutationsBasic_io_in_43_Im),
    .io_in_44_Re(PermutationsBasic_io_in_44_Re),
    .io_in_44_Im(PermutationsBasic_io_in_44_Im),
    .io_in_45_Re(PermutationsBasic_io_in_45_Re),
    .io_in_45_Im(PermutationsBasic_io_in_45_Im),
    .io_in_46_Re(PermutationsBasic_io_in_46_Re),
    .io_in_46_Im(PermutationsBasic_io_in_46_Im),
    .io_in_47_Re(PermutationsBasic_io_in_47_Re),
    .io_in_47_Im(PermutationsBasic_io_in_47_Im),
    .io_in_48_Re(PermutationsBasic_io_in_48_Re),
    .io_in_48_Im(PermutationsBasic_io_in_48_Im),
    .io_in_49_Re(PermutationsBasic_io_in_49_Re),
    .io_in_49_Im(PermutationsBasic_io_in_49_Im),
    .io_in_50_Re(PermutationsBasic_io_in_50_Re),
    .io_in_50_Im(PermutationsBasic_io_in_50_Im),
    .io_in_51_Re(PermutationsBasic_io_in_51_Re),
    .io_in_51_Im(PermutationsBasic_io_in_51_Im),
    .io_in_52_Re(PermutationsBasic_io_in_52_Re),
    .io_in_52_Im(PermutationsBasic_io_in_52_Im),
    .io_in_53_Re(PermutationsBasic_io_in_53_Re),
    .io_in_53_Im(PermutationsBasic_io_in_53_Im),
    .io_in_54_Re(PermutationsBasic_io_in_54_Re),
    .io_in_54_Im(PermutationsBasic_io_in_54_Im),
    .io_in_55_Re(PermutationsBasic_io_in_55_Re),
    .io_in_55_Im(PermutationsBasic_io_in_55_Im),
    .io_in_56_Re(PermutationsBasic_io_in_56_Re),
    .io_in_56_Im(PermutationsBasic_io_in_56_Im),
    .io_in_57_Re(PermutationsBasic_io_in_57_Re),
    .io_in_57_Im(PermutationsBasic_io_in_57_Im),
    .io_in_58_Re(PermutationsBasic_io_in_58_Re),
    .io_in_58_Im(PermutationsBasic_io_in_58_Im),
    .io_in_59_Re(PermutationsBasic_io_in_59_Re),
    .io_in_59_Im(PermutationsBasic_io_in_59_Im),
    .io_in_60_Re(PermutationsBasic_io_in_60_Re),
    .io_in_60_Im(PermutationsBasic_io_in_60_Im),
    .io_in_61_Re(PermutationsBasic_io_in_61_Re),
    .io_in_61_Im(PermutationsBasic_io_in_61_Im),
    .io_in_62_Re(PermutationsBasic_io_in_62_Re),
    .io_in_62_Im(PermutationsBasic_io_in_62_Im),
    .io_in_63_Re(PermutationsBasic_io_in_63_Re),
    .io_in_63_Im(PermutationsBasic_io_in_63_Im),
    .io_in_64_Re(PermutationsBasic_io_in_64_Re),
    .io_in_64_Im(PermutationsBasic_io_in_64_Im),
    .io_in_65_Re(PermutationsBasic_io_in_65_Re),
    .io_in_65_Im(PermutationsBasic_io_in_65_Im),
    .io_in_66_Re(PermutationsBasic_io_in_66_Re),
    .io_in_66_Im(PermutationsBasic_io_in_66_Im),
    .io_in_67_Re(PermutationsBasic_io_in_67_Re),
    .io_in_67_Im(PermutationsBasic_io_in_67_Im),
    .io_in_68_Re(PermutationsBasic_io_in_68_Re),
    .io_in_68_Im(PermutationsBasic_io_in_68_Im),
    .io_in_69_Re(PermutationsBasic_io_in_69_Re),
    .io_in_69_Im(PermutationsBasic_io_in_69_Im),
    .io_in_70_Re(PermutationsBasic_io_in_70_Re),
    .io_in_70_Im(PermutationsBasic_io_in_70_Im),
    .io_in_71_Re(PermutationsBasic_io_in_71_Re),
    .io_in_71_Im(PermutationsBasic_io_in_71_Im),
    .io_in_72_Re(PermutationsBasic_io_in_72_Re),
    .io_in_72_Im(PermutationsBasic_io_in_72_Im),
    .io_in_73_Re(PermutationsBasic_io_in_73_Re),
    .io_in_73_Im(PermutationsBasic_io_in_73_Im),
    .io_in_74_Re(PermutationsBasic_io_in_74_Re),
    .io_in_74_Im(PermutationsBasic_io_in_74_Im),
    .io_in_75_Re(PermutationsBasic_io_in_75_Re),
    .io_in_75_Im(PermutationsBasic_io_in_75_Im),
    .io_in_76_Re(PermutationsBasic_io_in_76_Re),
    .io_in_76_Im(PermutationsBasic_io_in_76_Im),
    .io_in_77_Re(PermutationsBasic_io_in_77_Re),
    .io_in_77_Im(PermutationsBasic_io_in_77_Im),
    .io_in_78_Re(PermutationsBasic_io_in_78_Re),
    .io_in_78_Im(PermutationsBasic_io_in_78_Im),
    .io_in_79_Re(PermutationsBasic_io_in_79_Re),
    .io_in_79_Im(PermutationsBasic_io_in_79_Im),
    .io_in_80_Re(PermutationsBasic_io_in_80_Re),
    .io_in_80_Im(PermutationsBasic_io_in_80_Im),
    .io_in_81_Re(PermutationsBasic_io_in_81_Re),
    .io_in_81_Im(PermutationsBasic_io_in_81_Im),
    .io_in_82_Re(PermutationsBasic_io_in_82_Re),
    .io_in_82_Im(PermutationsBasic_io_in_82_Im),
    .io_in_83_Re(PermutationsBasic_io_in_83_Re),
    .io_in_83_Im(PermutationsBasic_io_in_83_Im),
    .io_in_84_Re(PermutationsBasic_io_in_84_Re),
    .io_in_84_Im(PermutationsBasic_io_in_84_Im),
    .io_in_85_Re(PermutationsBasic_io_in_85_Re),
    .io_in_85_Im(PermutationsBasic_io_in_85_Im),
    .io_in_86_Re(PermutationsBasic_io_in_86_Re),
    .io_in_86_Im(PermutationsBasic_io_in_86_Im),
    .io_in_87_Re(PermutationsBasic_io_in_87_Re),
    .io_in_87_Im(PermutationsBasic_io_in_87_Im),
    .io_in_88_Re(PermutationsBasic_io_in_88_Re),
    .io_in_88_Im(PermutationsBasic_io_in_88_Im),
    .io_in_89_Re(PermutationsBasic_io_in_89_Re),
    .io_in_89_Im(PermutationsBasic_io_in_89_Im),
    .io_in_90_Re(PermutationsBasic_io_in_90_Re),
    .io_in_90_Im(PermutationsBasic_io_in_90_Im),
    .io_in_91_Re(PermutationsBasic_io_in_91_Re),
    .io_in_91_Im(PermutationsBasic_io_in_91_Im),
    .io_in_92_Re(PermutationsBasic_io_in_92_Re),
    .io_in_92_Im(PermutationsBasic_io_in_92_Im),
    .io_in_93_Re(PermutationsBasic_io_in_93_Re),
    .io_in_93_Im(PermutationsBasic_io_in_93_Im),
    .io_in_94_Re(PermutationsBasic_io_in_94_Re),
    .io_in_94_Im(PermutationsBasic_io_in_94_Im),
    .io_in_95_Re(PermutationsBasic_io_in_95_Re),
    .io_in_95_Im(PermutationsBasic_io_in_95_Im),
    .io_out_0_Re(PermutationsBasic_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_io_out_31_Im),
    .io_out_32_Re(PermutationsBasic_io_out_32_Re),
    .io_out_32_Im(PermutationsBasic_io_out_32_Im),
    .io_out_33_Re(PermutationsBasic_io_out_33_Re),
    .io_out_33_Im(PermutationsBasic_io_out_33_Im),
    .io_out_34_Re(PermutationsBasic_io_out_34_Re),
    .io_out_34_Im(PermutationsBasic_io_out_34_Im),
    .io_out_35_Re(PermutationsBasic_io_out_35_Re),
    .io_out_35_Im(PermutationsBasic_io_out_35_Im),
    .io_out_36_Re(PermutationsBasic_io_out_36_Re),
    .io_out_36_Im(PermutationsBasic_io_out_36_Im),
    .io_out_37_Re(PermutationsBasic_io_out_37_Re),
    .io_out_37_Im(PermutationsBasic_io_out_37_Im),
    .io_out_38_Re(PermutationsBasic_io_out_38_Re),
    .io_out_38_Im(PermutationsBasic_io_out_38_Im),
    .io_out_39_Re(PermutationsBasic_io_out_39_Re),
    .io_out_39_Im(PermutationsBasic_io_out_39_Im),
    .io_out_40_Re(PermutationsBasic_io_out_40_Re),
    .io_out_40_Im(PermutationsBasic_io_out_40_Im),
    .io_out_41_Re(PermutationsBasic_io_out_41_Re),
    .io_out_41_Im(PermutationsBasic_io_out_41_Im),
    .io_out_42_Re(PermutationsBasic_io_out_42_Re),
    .io_out_42_Im(PermutationsBasic_io_out_42_Im),
    .io_out_43_Re(PermutationsBasic_io_out_43_Re),
    .io_out_43_Im(PermutationsBasic_io_out_43_Im),
    .io_out_44_Re(PermutationsBasic_io_out_44_Re),
    .io_out_44_Im(PermutationsBasic_io_out_44_Im),
    .io_out_45_Re(PermutationsBasic_io_out_45_Re),
    .io_out_45_Im(PermutationsBasic_io_out_45_Im),
    .io_out_46_Re(PermutationsBasic_io_out_46_Re),
    .io_out_46_Im(PermutationsBasic_io_out_46_Im),
    .io_out_47_Re(PermutationsBasic_io_out_47_Re),
    .io_out_47_Im(PermutationsBasic_io_out_47_Im),
    .io_out_48_Re(PermutationsBasic_io_out_48_Re),
    .io_out_48_Im(PermutationsBasic_io_out_48_Im),
    .io_out_49_Re(PermutationsBasic_io_out_49_Re),
    .io_out_49_Im(PermutationsBasic_io_out_49_Im),
    .io_out_50_Re(PermutationsBasic_io_out_50_Re),
    .io_out_50_Im(PermutationsBasic_io_out_50_Im),
    .io_out_51_Re(PermutationsBasic_io_out_51_Re),
    .io_out_51_Im(PermutationsBasic_io_out_51_Im),
    .io_out_52_Re(PermutationsBasic_io_out_52_Re),
    .io_out_52_Im(PermutationsBasic_io_out_52_Im),
    .io_out_53_Re(PermutationsBasic_io_out_53_Re),
    .io_out_53_Im(PermutationsBasic_io_out_53_Im),
    .io_out_54_Re(PermutationsBasic_io_out_54_Re),
    .io_out_54_Im(PermutationsBasic_io_out_54_Im),
    .io_out_55_Re(PermutationsBasic_io_out_55_Re),
    .io_out_55_Im(PermutationsBasic_io_out_55_Im),
    .io_out_56_Re(PermutationsBasic_io_out_56_Re),
    .io_out_56_Im(PermutationsBasic_io_out_56_Im),
    .io_out_57_Re(PermutationsBasic_io_out_57_Re),
    .io_out_57_Im(PermutationsBasic_io_out_57_Im),
    .io_out_58_Re(PermutationsBasic_io_out_58_Re),
    .io_out_58_Im(PermutationsBasic_io_out_58_Im),
    .io_out_59_Re(PermutationsBasic_io_out_59_Re),
    .io_out_59_Im(PermutationsBasic_io_out_59_Im),
    .io_out_60_Re(PermutationsBasic_io_out_60_Re),
    .io_out_60_Im(PermutationsBasic_io_out_60_Im),
    .io_out_61_Re(PermutationsBasic_io_out_61_Re),
    .io_out_61_Im(PermutationsBasic_io_out_61_Im),
    .io_out_62_Re(PermutationsBasic_io_out_62_Re),
    .io_out_62_Im(PermutationsBasic_io_out_62_Im),
    .io_out_63_Re(PermutationsBasic_io_out_63_Re),
    .io_out_63_Im(PermutationsBasic_io_out_63_Im),
    .io_out_64_Re(PermutationsBasic_io_out_64_Re),
    .io_out_64_Im(PermutationsBasic_io_out_64_Im),
    .io_out_65_Re(PermutationsBasic_io_out_65_Re),
    .io_out_65_Im(PermutationsBasic_io_out_65_Im),
    .io_out_66_Re(PermutationsBasic_io_out_66_Re),
    .io_out_66_Im(PermutationsBasic_io_out_66_Im),
    .io_out_67_Re(PermutationsBasic_io_out_67_Re),
    .io_out_67_Im(PermutationsBasic_io_out_67_Im),
    .io_out_68_Re(PermutationsBasic_io_out_68_Re),
    .io_out_68_Im(PermutationsBasic_io_out_68_Im),
    .io_out_69_Re(PermutationsBasic_io_out_69_Re),
    .io_out_69_Im(PermutationsBasic_io_out_69_Im),
    .io_out_70_Re(PermutationsBasic_io_out_70_Re),
    .io_out_70_Im(PermutationsBasic_io_out_70_Im),
    .io_out_71_Re(PermutationsBasic_io_out_71_Re),
    .io_out_71_Im(PermutationsBasic_io_out_71_Im),
    .io_out_72_Re(PermutationsBasic_io_out_72_Re),
    .io_out_72_Im(PermutationsBasic_io_out_72_Im),
    .io_out_73_Re(PermutationsBasic_io_out_73_Re),
    .io_out_73_Im(PermutationsBasic_io_out_73_Im),
    .io_out_74_Re(PermutationsBasic_io_out_74_Re),
    .io_out_74_Im(PermutationsBasic_io_out_74_Im),
    .io_out_75_Re(PermutationsBasic_io_out_75_Re),
    .io_out_75_Im(PermutationsBasic_io_out_75_Im),
    .io_out_76_Re(PermutationsBasic_io_out_76_Re),
    .io_out_76_Im(PermutationsBasic_io_out_76_Im),
    .io_out_77_Re(PermutationsBasic_io_out_77_Re),
    .io_out_77_Im(PermutationsBasic_io_out_77_Im),
    .io_out_78_Re(PermutationsBasic_io_out_78_Re),
    .io_out_78_Im(PermutationsBasic_io_out_78_Im),
    .io_out_79_Re(PermutationsBasic_io_out_79_Re),
    .io_out_79_Im(PermutationsBasic_io_out_79_Im),
    .io_out_80_Re(PermutationsBasic_io_out_80_Re),
    .io_out_80_Im(PermutationsBasic_io_out_80_Im),
    .io_out_81_Re(PermutationsBasic_io_out_81_Re),
    .io_out_81_Im(PermutationsBasic_io_out_81_Im),
    .io_out_82_Re(PermutationsBasic_io_out_82_Re),
    .io_out_82_Im(PermutationsBasic_io_out_82_Im),
    .io_out_83_Re(PermutationsBasic_io_out_83_Re),
    .io_out_83_Im(PermutationsBasic_io_out_83_Im),
    .io_out_84_Re(PermutationsBasic_io_out_84_Re),
    .io_out_84_Im(PermutationsBasic_io_out_84_Im),
    .io_out_85_Re(PermutationsBasic_io_out_85_Re),
    .io_out_85_Im(PermutationsBasic_io_out_85_Im),
    .io_out_86_Re(PermutationsBasic_io_out_86_Re),
    .io_out_86_Im(PermutationsBasic_io_out_86_Im),
    .io_out_87_Re(PermutationsBasic_io_out_87_Re),
    .io_out_87_Im(PermutationsBasic_io_out_87_Im),
    .io_out_88_Re(PermutationsBasic_io_out_88_Re),
    .io_out_88_Im(PermutationsBasic_io_out_88_Im),
    .io_out_89_Re(PermutationsBasic_io_out_89_Re),
    .io_out_89_Im(PermutationsBasic_io_out_89_Im),
    .io_out_90_Re(PermutationsBasic_io_out_90_Re),
    .io_out_90_Im(PermutationsBasic_io_out_90_Im),
    .io_out_91_Re(PermutationsBasic_io_out_91_Re),
    .io_out_91_Im(PermutationsBasic_io_out_91_Im),
    .io_out_92_Re(PermutationsBasic_io_out_92_Re),
    .io_out_92_Im(PermutationsBasic_io_out_92_Im),
    .io_out_93_Re(PermutationsBasic_io_out_93_Re),
    .io_out_93_Im(PermutationsBasic_io_out_93_Im),
    .io_out_94_Re(PermutationsBasic_io_out_94_Re),
    .io_out_94_Im(PermutationsBasic_io_out_94_Im),
    .io_out_95_Re(PermutationsBasic_io_out_95_Re),
    .io_out_95_Im(PermutationsBasic_io_out_95_Im)
  );
  PermutationsBasic_83 PermutationsBasic_1 ( // @[FFTDesigns.scala 3447:27]
    .io_in_0_Re(PermutationsBasic_1_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_1_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_1_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_1_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_1_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_1_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_1_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_1_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_1_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_1_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_1_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_1_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_1_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_1_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_1_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_1_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_1_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_1_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_1_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_1_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_1_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_1_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_1_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_1_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_1_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_1_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_1_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_1_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_1_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_1_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_1_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_1_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_1_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_1_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_1_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_1_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_1_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_1_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_1_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_1_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_1_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_1_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_1_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_1_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_1_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_1_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_1_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_1_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_1_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_1_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_1_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_1_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_1_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_1_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_1_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_1_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_1_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_1_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_1_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_1_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_1_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_1_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_1_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_1_io_in_31_Im),
    .io_in_32_Re(PermutationsBasic_1_io_in_32_Re),
    .io_in_32_Im(PermutationsBasic_1_io_in_32_Im),
    .io_in_33_Re(PermutationsBasic_1_io_in_33_Re),
    .io_in_33_Im(PermutationsBasic_1_io_in_33_Im),
    .io_in_34_Re(PermutationsBasic_1_io_in_34_Re),
    .io_in_34_Im(PermutationsBasic_1_io_in_34_Im),
    .io_in_35_Re(PermutationsBasic_1_io_in_35_Re),
    .io_in_35_Im(PermutationsBasic_1_io_in_35_Im),
    .io_in_36_Re(PermutationsBasic_1_io_in_36_Re),
    .io_in_36_Im(PermutationsBasic_1_io_in_36_Im),
    .io_in_37_Re(PermutationsBasic_1_io_in_37_Re),
    .io_in_37_Im(PermutationsBasic_1_io_in_37_Im),
    .io_in_38_Re(PermutationsBasic_1_io_in_38_Re),
    .io_in_38_Im(PermutationsBasic_1_io_in_38_Im),
    .io_in_39_Re(PermutationsBasic_1_io_in_39_Re),
    .io_in_39_Im(PermutationsBasic_1_io_in_39_Im),
    .io_in_40_Re(PermutationsBasic_1_io_in_40_Re),
    .io_in_40_Im(PermutationsBasic_1_io_in_40_Im),
    .io_in_41_Re(PermutationsBasic_1_io_in_41_Re),
    .io_in_41_Im(PermutationsBasic_1_io_in_41_Im),
    .io_in_42_Re(PermutationsBasic_1_io_in_42_Re),
    .io_in_42_Im(PermutationsBasic_1_io_in_42_Im),
    .io_in_43_Re(PermutationsBasic_1_io_in_43_Re),
    .io_in_43_Im(PermutationsBasic_1_io_in_43_Im),
    .io_in_44_Re(PermutationsBasic_1_io_in_44_Re),
    .io_in_44_Im(PermutationsBasic_1_io_in_44_Im),
    .io_in_45_Re(PermutationsBasic_1_io_in_45_Re),
    .io_in_45_Im(PermutationsBasic_1_io_in_45_Im),
    .io_in_46_Re(PermutationsBasic_1_io_in_46_Re),
    .io_in_46_Im(PermutationsBasic_1_io_in_46_Im),
    .io_in_47_Re(PermutationsBasic_1_io_in_47_Re),
    .io_in_47_Im(PermutationsBasic_1_io_in_47_Im),
    .io_in_48_Re(PermutationsBasic_1_io_in_48_Re),
    .io_in_48_Im(PermutationsBasic_1_io_in_48_Im),
    .io_in_49_Re(PermutationsBasic_1_io_in_49_Re),
    .io_in_49_Im(PermutationsBasic_1_io_in_49_Im),
    .io_in_50_Re(PermutationsBasic_1_io_in_50_Re),
    .io_in_50_Im(PermutationsBasic_1_io_in_50_Im),
    .io_in_51_Re(PermutationsBasic_1_io_in_51_Re),
    .io_in_51_Im(PermutationsBasic_1_io_in_51_Im),
    .io_in_52_Re(PermutationsBasic_1_io_in_52_Re),
    .io_in_52_Im(PermutationsBasic_1_io_in_52_Im),
    .io_in_53_Re(PermutationsBasic_1_io_in_53_Re),
    .io_in_53_Im(PermutationsBasic_1_io_in_53_Im),
    .io_in_54_Re(PermutationsBasic_1_io_in_54_Re),
    .io_in_54_Im(PermutationsBasic_1_io_in_54_Im),
    .io_in_55_Re(PermutationsBasic_1_io_in_55_Re),
    .io_in_55_Im(PermutationsBasic_1_io_in_55_Im),
    .io_in_56_Re(PermutationsBasic_1_io_in_56_Re),
    .io_in_56_Im(PermutationsBasic_1_io_in_56_Im),
    .io_in_57_Re(PermutationsBasic_1_io_in_57_Re),
    .io_in_57_Im(PermutationsBasic_1_io_in_57_Im),
    .io_in_58_Re(PermutationsBasic_1_io_in_58_Re),
    .io_in_58_Im(PermutationsBasic_1_io_in_58_Im),
    .io_in_59_Re(PermutationsBasic_1_io_in_59_Re),
    .io_in_59_Im(PermutationsBasic_1_io_in_59_Im),
    .io_in_60_Re(PermutationsBasic_1_io_in_60_Re),
    .io_in_60_Im(PermutationsBasic_1_io_in_60_Im),
    .io_in_61_Re(PermutationsBasic_1_io_in_61_Re),
    .io_in_61_Im(PermutationsBasic_1_io_in_61_Im),
    .io_in_62_Re(PermutationsBasic_1_io_in_62_Re),
    .io_in_62_Im(PermutationsBasic_1_io_in_62_Im),
    .io_in_63_Re(PermutationsBasic_1_io_in_63_Re),
    .io_in_63_Im(PermutationsBasic_1_io_in_63_Im),
    .io_in_64_Re(PermutationsBasic_1_io_in_64_Re),
    .io_in_64_Im(PermutationsBasic_1_io_in_64_Im),
    .io_in_65_Re(PermutationsBasic_1_io_in_65_Re),
    .io_in_65_Im(PermutationsBasic_1_io_in_65_Im),
    .io_in_66_Re(PermutationsBasic_1_io_in_66_Re),
    .io_in_66_Im(PermutationsBasic_1_io_in_66_Im),
    .io_in_67_Re(PermutationsBasic_1_io_in_67_Re),
    .io_in_67_Im(PermutationsBasic_1_io_in_67_Im),
    .io_in_68_Re(PermutationsBasic_1_io_in_68_Re),
    .io_in_68_Im(PermutationsBasic_1_io_in_68_Im),
    .io_in_69_Re(PermutationsBasic_1_io_in_69_Re),
    .io_in_69_Im(PermutationsBasic_1_io_in_69_Im),
    .io_in_70_Re(PermutationsBasic_1_io_in_70_Re),
    .io_in_70_Im(PermutationsBasic_1_io_in_70_Im),
    .io_in_71_Re(PermutationsBasic_1_io_in_71_Re),
    .io_in_71_Im(PermutationsBasic_1_io_in_71_Im),
    .io_in_72_Re(PermutationsBasic_1_io_in_72_Re),
    .io_in_72_Im(PermutationsBasic_1_io_in_72_Im),
    .io_in_73_Re(PermutationsBasic_1_io_in_73_Re),
    .io_in_73_Im(PermutationsBasic_1_io_in_73_Im),
    .io_in_74_Re(PermutationsBasic_1_io_in_74_Re),
    .io_in_74_Im(PermutationsBasic_1_io_in_74_Im),
    .io_in_75_Re(PermutationsBasic_1_io_in_75_Re),
    .io_in_75_Im(PermutationsBasic_1_io_in_75_Im),
    .io_in_76_Re(PermutationsBasic_1_io_in_76_Re),
    .io_in_76_Im(PermutationsBasic_1_io_in_76_Im),
    .io_in_77_Re(PermutationsBasic_1_io_in_77_Re),
    .io_in_77_Im(PermutationsBasic_1_io_in_77_Im),
    .io_in_78_Re(PermutationsBasic_1_io_in_78_Re),
    .io_in_78_Im(PermutationsBasic_1_io_in_78_Im),
    .io_in_79_Re(PermutationsBasic_1_io_in_79_Re),
    .io_in_79_Im(PermutationsBasic_1_io_in_79_Im),
    .io_in_80_Re(PermutationsBasic_1_io_in_80_Re),
    .io_in_80_Im(PermutationsBasic_1_io_in_80_Im),
    .io_in_81_Re(PermutationsBasic_1_io_in_81_Re),
    .io_in_81_Im(PermutationsBasic_1_io_in_81_Im),
    .io_in_82_Re(PermutationsBasic_1_io_in_82_Re),
    .io_in_82_Im(PermutationsBasic_1_io_in_82_Im),
    .io_in_83_Re(PermutationsBasic_1_io_in_83_Re),
    .io_in_83_Im(PermutationsBasic_1_io_in_83_Im),
    .io_in_84_Re(PermutationsBasic_1_io_in_84_Re),
    .io_in_84_Im(PermutationsBasic_1_io_in_84_Im),
    .io_in_85_Re(PermutationsBasic_1_io_in_85_Re),
    .io_in_85_Im(PermutationsBasic_1_io_in_85_Im),
    .io_in_86_Re(PermutationsBasic_1_io_in_86_Re),
    .io_in_86_Im(PermutationsBasic_1_io_in_86_Im),
    .io_in_87_Re(PermutationsBasic_1_io_in_87_Re),
    .io_in_87_Im(PermutationsBasic_1_io_in_87_Im),
    .io_in_88_Re(PermutationsBasic_1_io_in_88_Re),
    .io_in_88_Im(PermutationsBasic_1_io_in_88_Im),
    .io_in_89_Re(PermutationsBasic_1_io_in_89_Re),
    .io_in_89_Im(PermutationsBasic_1_io_in_89_Im),
    .io_in_90_Re(PermutationsBasic_1_io_in_90_Re),
    .io_in_90_Im(PermutationsBasic_1_io_in_90_Im),
    .io_in_91_Re(PermutationsBasic_1_io_in_91_Re),
    .io_in_91_Im(PermutationsBasic_1_io_in_91_Im),
    .io_in_92_Re(PermutationsBasic_1_io_in_92_Re),
    .io_in_92_Im(PermutationsBasic_1_io_in_92_Im),
    .io_in_93_Re(PermutationsBasic_1_io_in_93_Re),
    .io_in_93_Im(PermutationsBasic_1_io_in_93_Im),
    .io_in_94_Re(PermutationsBasic_1_io_in_94_Re),
    .io_in_94_Im(PermutationsBasic_1_io_in_94_Im),
    .io_in_95_Re(PermutationsBasic_1_io_in_95_Re),
    .io_in_95_Im(PermutationsBasic_1_io_in_95_Im),
    .io_out_0_Re(PermutationsBasic_1_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_1_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_1_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_1_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_1_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_1_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_1_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_1_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_1_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_1_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_1_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_1_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_1_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_1_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_1_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_1_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_1_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_1_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_1_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_1_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_1_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_1_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_1_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_1_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_1_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_1_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_1_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_1_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_1_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_1_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_1_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_1_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_1_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_1_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_1_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_1_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_1_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_1_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_1_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_1_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_1_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_1_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_1_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_1_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_1_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_1_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_1_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_1_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_1_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_1_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_1_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_1_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_1_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_1_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_1_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_1_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_1_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_1_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_1_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_1_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_1_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_1_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_1_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_1_io_out_31_Im),
    .io_out_32_Re(PermutationsBasic_1_io_out_32_Re),
    .io_out_32_Im(PermutationsBasic_1_io_out_32_Im),
    .io_out_33_Re(PermutationsBasic_1_io_out_33_Re),
    .io_out_33_Im(PermutationsBasic_1_io_out_33_Im),
    .io_out_34_Re(PermutationsBasic_1_io_out_34_Re),
    .io_out_34_Im(PermutationsBasic_1_io_out_34_Im),
    .io_out_35_Re(PermutationsBasic_1_io_out_35_Re),
    .io_out_35_Im(PermutationsBasic_1_io_out_35_Im),
    .io_out_36_Re(PermutationsBasic_1_io_out_36_Re),
    .io_out_36_Im(PermutationsBasic_1_io_out_36_Im),
    .io_out_37_Re(PermutationsBasic_1_io_out_37_Re),
    .io_out_37_Im(PermutationsBasic_1_io_out_37_Im),
    .io_out_38_Re(PermutationsBasic_1_io_out_38_Re),
    .io_out_38_Im(PermutationsBasic_1_io_out_38_Im),
    .io_out_39_Re(PermutationsBasic_1_io_out_39_Re),
    .io_out_39_Im(PermutationsBasic_1_io_out_39_Im),
    .io_out_40_Re(PermutationsBasic_1_io_out_40_Re),
    .io_out_40_Im(PermutationsBasic_1_io_out_40_Im),
    .io_out_41_Re(PermutationsBasic_1_io_out_41_Re),
    .io_out_41_Im(PermutationsBasic_1_io_out_41_Im),
    .io_out_42_Re(PermutationsBasic_1_io_out_42_Re),
    .io_out_42_Im(PermutationsBasic_1_io_out_42_Im),
    .io_out_43_Re(PermutationsBasic_1_io_out_43_Re),
    .io_out_43_Im(PermutationsBasic_1_io_out_43_Im),
    .io_out_44_Re(PermutationsBasic_1_io_out_44_Re),
    .io_out_44_Im(PermutationsBasic_1_io_out_44_Im),
    .io_out_45_Re(PermutationsBasic_1_io_out_45_Re),
    .io_out_45_Im(PermutationsBasic_1_io_out_45_Im),
    .io_out_46_Re(PermutationsBasic_1_io_out_46_Re),
    .io_out_46_Im(PermutationsBasic_1_io_out_46_Im),
    .io_out_47_Re(PermutationsBasic_1_io_out_47_Re),
    .io_out_47_Im(PermutationsBasic_1_io_out_47_Im),
    .io_out_48_Re(PermutationsBasic_1_io_out_48_Re),
    .io_out_48_Im(PermutationsBasic_1_io_out_48_Im),
    .io_out_49_Re(PermutationsBasic_1_io_out_49_Re),
    .io_out_49_Im(PermutationsBasic_1_io_out_49_Im),
    .io_out_50_Re(PermutationsBasic_1_io_out_50_Re),
    .io_out_50_Im(PermutationsBasic_1_io_out_50_Im),
    .io_out_51_Re(PermutationsBasic_1_io_out_51_Re),
    .io_out_51_Im(PermutationsBasic_1_io_out_51_Im),
    .io_out_52_Re(PermutationsBasic_1_io_out_52_Re),
    .io_out_52_Im(PermutationsBasic_1_io_out_52_Im),
    .io_out_53_Re(PermutationsBasic_1_io_out_53_Re),
    .io_out_53_Im(PermutationsBasic_1_io_out_53_Im),
    .io_out_54_Re(PermutationsBasic_1_io_out_54_Re),
    .io_out_54_Im(PermutationsBasic_1_io_out_54_Im),
    .io_out_55_Re(PermutationsBasic_1_io_out_55_Re),
    .io_out_55_Im(PermutationsBasic_1_io_out_55_Im),
    .io_out_56_Re(PermutationsBasic_1_io_out_56_Re),
    .io_out_56_Im(PermutationsBasic_1_io_out_56_Im),
    .io_out_57_Re(PermutationsBasic_1_io_out_57_Re),
    .io_out_57_Im(PermutationsBasic_1_io_out_57_Im),
    .io_out_58_Re(PermutationsBasic_1_io_out_58_Re),
    .io_out_58_Im(PermutationsBasic_1_io_out_58_Im),
    .io_out_59_Re(PermutationsBasic_1_io_out_59_Re),
    .io_out_59_Im(PermutationsBasic_1_io_out_59_Im),
    .io_out_60_Re(PermutationsBasic_1_io_out_60_Re),
    .io_out_60_Im(PermutationsBasic_1_io_out_60_Im),
    .io_out_61_Re(PermutationsBasic_1_io_out_61_Re),
    .io_out_61_Im(PermutationsBasic_1_io_out_61_Im),
    .io_out_62_Re(PermutationsBasic_1_io_out_62_Re),
    .io_out_62_Im(PermutationsBasic_1_io_out_62_Im),
    .io_out_63_Re(PermutationsBasic_1_io_out_63_Re),
    .io_out_63_Im(PermutationsBasic_1_io_out_63_Im),
    .io_out_64_Re(PermutationsBasic_1_io_out_64_Re),
    .io_out_64_Im(PermutationsBasic_1_io_out_64_Im),
    .io_out_65_Re(PermutationsBasic_1_io_out_65_Re),
    .io_out_65_Im(PermutationsBasic_1_io_out_65_Im),
    .io_out_66_Re(PermutationsBasic_1_io_out_66_Re),
    .io_out_66_Im(PermutationsBasic_1_io_out_66_Im),
    .io_out_67_Re(PermutationsBasic_1_io_out_67_Re),
    .io_out_67_Im(PermutationsBasic_1_io_out_67_Im),
    .io_out_68_Re(PermutationsBasic_1_io_out_68_Re),
    .io_out_68_Im(PermutationsBasic_1_io_out_68_Im),
    .io_out_69_Re(PermutationsBasic_1_io_out_69_Re),
    .io_out_69_Im(PermutationsBasic_1_io_out_69_Im),
    .io_out_70_Re(PermutationsBasic_1_io_out_70_Re),
    .io_out_70_Im(PermutationsBasic_1_io_out_70_Im),
    .io_out_71_Re(PermutationsBasic_1_io_out_71_Re),
    .io_out_71_Im(PermutationsBasic_1_io_out_71_Im),
    .io_out_72_Re(PermutationsBasic_1_io_out_72_Re),
    .io_out_72_Im(PermutationsBasic_1_io_out_72_Im),
    .io_out_73_Re(PermutationsBasic_1_io_out_73_Re),
    .io_out_73_Im(PermutationsBasic_1_io_out_73_Im),
    .io_out_74_Re(PermutationsBasic_1_io_out_74_Re),
    .io_out_74_Im(PermutationsBasic_1_io_out_74_Im),
    .io_out_75_Re(PermutationsBasic_1_io_out_75_Re),
    .io_out_75_Im(PermutationsBasic_1_io_out_75_Im),
    .io_out_76_Re(PermutationsBasic_1_io_out_76_Re),
    .io_out_76_Im(PermutationsBasic_1_io_out_76_Im),
    .io_out_77_Re(PermutationsBasic_1_io_out_77_Re),
    .io_out_77_Im(PermutationsBasic_1_io_out_77_Im),
    .io_out_78_Re(PermutationsBasic_1_io_out_78_Re),
    .io_out_78_Im(PermutationsBasic_1_io_out_78_Im),
    .io_out_79_Re(PermutationsBasic_1_io_out_79_Re),
    .io_out_79_Im(PermutationsBasic_1_io_out_79_Im),
    .io_out_80_Re(PermutationsBasic_1_io_out_80_Re),
    .io_out_80_Im(PermutationsBasic_1_io_out_80_Im),
    .io_out_81_Re(PermutationsBasic_1_io_out_81_Re),
    .io_out_81_Im(PermutationsBasic_1_io_out_81_Im),
    .io_out_82_Re(PermutationsBasic_1_io_out_82_Re),
    .io_out_82_Im(PermutationsBasic_1_io_out_82_Im),
    .io_out_83_Re(PermutationsBasic_1_io_out_83_Re),
    .io_out_83_Im(PermutationsBasic_1_io_out_83_Im),
    .io_out_84_Re(PermutationsBasic_1_io_out_84_Re),
    .io_out_84_Im(PermutationsBasic_1_io_out_84_Im),
    .io_out_85_Re(PermutationsBasic_1_io_out_85_Re),
    .io_out_85_Im(PermutationsBasic_1_io_out_85_Im),
    .io_out_86_Re(PermutationsBasic_1_io_out_86_Re),
    .io_out_86_Im(PermutationsBasic_1_io_out_86_Im),
    .io_out_87_Re(PermutationsBasic_1_io_out_87_Re),
    .io_out_87_Im(PermutationsBasic_1_io_out_87_Im),
    .io_out_88_Re(PermutationsBasic_1_io_out_88_Re),
    .io_out_88_Im(PermutationsBasic_1_io_out_88_Im),
    .io_out_89_Re(PermutationsBasic_1_io_out_89_Re),
    .io_out_89_Im(PermutationsBasic_1_io_out_89_Im),
    .io_out_90_Re(PermutationsBasic_1_io_out_90_Re),
    .io_out_90_Im(PermutationsBasic_1_io_out_90_Im),
    .io_out_91_Re(PermutationsBasic_1_io_out_91_Re),
    .io_out_91_Im(PermutationsBasic_1_io_out_91_Im),
    .io_out_92_Re(PermutationsBasic_1_io_out_92_Re),
    .io_out_92_Im(PermutationsBasic_1_io_out_92_Im),
    .io_out_93_Re(PermutationsBasic_1_io_out_93_Re),
    .io_out_93_Im(PermutationsBasic_1_io_out_93_Im),
    .io_out_94_Re(PermutationsBasic_1_io_out_94_Re),
    .io_out_94_Im(PermutationsBasic_1_io_out_94_Im),
    .io_out_95_Re(PermutationsBasic_1_io_out_95_Re),
    .io_out_95_Im(PermutationsBasic_1_io_out_95_Im)
  );
  PermutationsBasic_82 PermutationsBasic_2 ( // @[FFTDesigns.scala 3450:27]
    .io_in_0_Re(PermutationsBasic_2_io_in_0_Re),
    .io_in_0_Im(PermutationsBasic_2_io_in_0_Im),
    .io_in_1_Re(PermutationsBasic_2_io_in_1_Re),
    .io_in_1_Im(PermutationsBasic_2_io_in_1_Im),
    .io_in_2_Re(PermutationsBasic_2_io_in_2_Re),
    .io_in_2_Im(PermutationsBasic_2_io_in_2_Im),
    .io_in_3_Re(PermutationsBasic_2_io_in_3_Re),
    .io_in_3_Im(PermutationsBasic_2_io_in_3_Im),
    .io_in_4_Re(PermutationsBasic_2_io_in_4_Re),
    .io_in_4_Im(PermutationsBasic_2_io_in_4_Im),
    .io_in_5_Re(PermutationsBasic_2_io_in_5_Re),
    .io_in_5_Im(PermutationsBasic_2_io_in_5_Im),
    .io_in_6_Re(PermutationsBasic_2_io_in_6_Re),
    .io_in_6_Im(PermutationsBasic_2_io_in_6_Im),
    .io_in_7_Re(PermutationsBasic_2_io_in_7_Re),
    .io_in_7_Im(PermutationsBasic_2_io_in_7_Im),
    .io_in_8_Re(PermutationsBasic_2_io_in_8_Re),
    .io_in_8_Im(PermutationsBasic_2_io_in_8_Im),
    .io_in_9_Re(PermutationsBasic_2_io_in_9_Re),
    .io_in_9_Im(PermutationsBasic_2_io_in_9_Im),
    .io_in_10_Re(PermutationsBasic_2_io_in_10_Re),
    .io_in_10_Im(PermutationsBasic_2_io_in_10_Im),
    .io_in_11_Re(PermutationsBasic_2_io_in_11_Re),
    .io_in_11_Im(PermutationsBasic_2_io_in_11_Im),
    .io_in_12_Re(PermutationsBasic_2_io_in_12_Re),
    .io_in_12_Im(PermutationsBasic_2_io_in_12_Im),
    .io_in_13_Re(PermutationsBasic_2_io_in_13_Re),
    .io_in_13_Im(PermutationsBasic_2_io_in_13_Im),
    .io_in_14_Re(PermutationsBasic_2_io_in_14_Re),
    .io_in_14_Im(PermutationsBasic_2_io_in_14_Im),
    .io_in_15_Re(PermutationsBasic_2_io_in_15_Re),
    .io_in_15_Im(PermutationsBasic_2_io_in_15_Im),
    .io_in_16_Re(PermutationsBasic_2_io_in_16_Re),
    .io_in_16_Im(PermutationsBasic_2_io_in_16_Im),
    .io_in_17_Re(PermutationsBasic_2_io_in_17_Re),
    .io_in_17_Im(PermutationsBasic_2_io_in_17_Im),
    .io_in_18_Re(PermutationsBasic_2_io_in_18_Re),
    .io_in_18_Im(PermutationsBasic_2_io_in_18_Im),
    .io_in_19_Re(PermutationsBasic_2_io_in_19_Re),
    .io_in_19_Im(PermutationsBasic_2_io_in_19_Im),
    .io_in_20_Re(PermutationsBasic_2_io_in_20_Re),
    .io_in_20_Im(PermutationsBasic_2_io_in_20_Im),
    .io_in_21_Re(PermutationsBasic_2_io_in_21_Re),
    .io_in_21_Im(PermutationsBasic_2_io_in_21_Im),
    .io_in_22_Re(PermutationsBasic_2_io_in_22_Re),
    .io_in_22_Im(PermutationsBasic_2_io_in_22_Im),
    .io_in_23_Re(PermutationsBasic_2_io_in_23_Re),
    .io_in_23_Im(PermutationsBasic_2_io_in_23_Im),
    .io_in_24_Re(PermutationsBasic_2_io_in_24_Re),
    .io_in_24_Im(PermutationsBasic_2_io_in_24_Im),
    .io_in_25_Re(PermutationsBasic_2_io_in_25_Re),
    .io_in_25_Im(PermutationsBasic_2_io_in_25_Im),
    .io_in_26_Re(PermutationsBasic_2_io_in_26_Re),
    .io_in_26_Im(PermutationsBasic_2_io_in_26_Im),
    .io_in_27_Re(PermutationsBasic_2_io_in_27_Re),
    .io_in_27_Im(PermutationsBasic_2_io_in_27_Im),
    .io_in_28_Re(PermutationsBasic_2_io_in_28_Re),
    .io_in_28_Im(PermutationsBasic_2_io_in_28_Im),
    .io_in_29_Re(PermutationsBasic_2_io_in_29_Re),
    .io_in_29_Im(PermutationsBasic_2_io_in_29_Im),
    .io_in_30_Re(PermutationsBasic_2_io_in_30_Re),
    .io_in_30_Im(PermutationsBasic_2_io_in_30_Im),
    .io_in_31_Re(PermutationsBasic_2_io_in_31_Re),
    .io_in_31_Im(PermutationsBasic_2_io_in_31_Im),
    .io_in_32_Re(PermutationsBasic_2_io_in_32_Re),
    .io_in_32_Im(PermutationsBasic_2_io_in_32_Im),
    .io_in_33_Re(PermutationsBasic_2_io_in_33_Re),
    .io_in_33_Im(PermutationsBasic_2_io_in_33_Im),
    .io_in_34_Re(PermutationsBasic_2_io_in_34_Re),
    .io_in_34_Im(PermutationsBasic_2_io_in_34_Im),
    .io_in_35_Re(PermutationsBasic_2_io_in_35_Re),
    .io_in_35_Im(PermutationsBasic_2_io_in_35_Im),
    .io_in_36_Re(PermutationsBasic_2_io_in_36_Re),
    .io_in_36_Im(PermutationsBasic_2_io_in_36_Im),
    .io_in_37_Re(PermutationsBasic_2_io_in_37_Re),
    .io_in_37_Im(PermutationsBasic_2_io_in_37_Im),
    .io_in_38_Re(PermutationsBasic_2_io_in_38_Re),
    .io_in_38_Im(PermutationsBasic_2_io_in_38_Im),
    .io_in_39_Re(PermutationsBasic_2_io_in_39_Re),
    .io_in_39_Im(PermutationsBasic_2_io_in_39_Im),
    .io_in_40_Re(PermutationsBasic_2_io_in_40_Re),
    .io_in_40_Im(PermutationsBasic_2_io_in_40_Im),
    .io_in_41_Re(PermutationsBasic_2_io_in_41_Re),
    .io_in_41_Im(PermutationsBasic_2_io_in_41_Im),
    .io_in_42_Re(PermutationsBasic_2_io_in_42_Re),
    .io_in_42_Im(PermutationsBasic_2_io_in_42_Im),
    .io_in_43_Re(PermutationsBasic_2_io_in_43_Re),
    .io_in_43_Im(PermutationsBasic_2_io_in_43_Im),
    .io_in_44_Re(PermutationsBasic_2_io_in_44_Re),
    .io_in_44_Im(PermutationsBasic_2_io_in_44_Im),
    .io_in_45_Re(PermutationsBasic_2_io_in_45_Re),
    .io_in_45_Im(PermutationsBasic_2_io_in_45_Im),
    .io_in_46_Re(PermutationsBasic_2_io_in_46_Re),
    .io_in_46_Im(PermutationsBasic_2_io_in_46_Im),
    .io_in_47_Re(PermutationsBasic_2_io_in_47_Re),
    .io_in_47_Im(PermutationsBasic_2_io_in_47_Im),
    .io_in_48_Re(PermutationsBasic_2_io_in_48_Re),
    .io_in_48_Im(PermutationsBasic_2_io_in_48_Im),
    .io_in_49_Re(PermutationsBasic_2_io_in_49_Re),
    .io_in_49_Im(PermutationsBasic_2_io_in_49_Im),
    .io_in_50_Re(PermutationsBasic_2_io_in_50_Re),
    .io_in_50_Im(PermutationsBasic_2_io_in_50_Im),
    .io_in_51_Re(PermutationsBasic_2_io_in_51_Re),
    .io_in_51_Im(PermutationsBasic_2_io_in_51_Im),
    .io_in_52_Re(PermutationsBasic_2_io_in_52_Re),
    .io_in_52_Im(PermutationsBasic_2_io_in_52_Im),
    .io_in_53_Re(PermutationsBasic_2_io_in_53_Re),
    .io_in_53_Im(PermutationsBasic_2_io_in_53_Im),
    .io_in_54_Re(PermutationsBasic_2_io_in_54_Re),
    .io_in_54_Im(PermutationsBasic_2_io_in_54_Im),
    .io_in_55_Re(PermutationsBasic_2_io_in_55_Re),
    .io_in_55_Im(PermutationsBasic_2_io_in_55_Im),
    .io_in_56_Re(PermutationsBasic_2_io_in_56_Re),
    .io_in_56_Im(PermutationsBasic_2_io_in_56_Im),
    .io_in_57_Re(PermutationsBasic_2_io_in_57_Re),
    .io_in_57_Im(PermutationsBasic_2_io_in_57_Im),
    .io_in_58_Re(PermutationsBasic_2_io_in_58_Re),
    .io_in_58_Im(PermutationsBasic_2_io_in_58_Im),
    .io_in_59_Re(PermutationsBasic_2_io_in_59_Re),
    .io_in_59_Im(PermutationsBasic_2_io_in_59_Im),
    .io_in_60_Re(PermutationsBasic_2_io_in_60_Re),
    .io_in_60_Im(PermutationsBasic_2_io_in_60_Im),
    .io_in_61_Re(PermutationsBasic_2_io_in_61_Re),
    .io_in_61_Im(PermutationsBasic_2_io_in_61_Im),
    .io_in_62_Re(PermutationsBasic_2_io_in_62_Re),
    .io_in_62_Im(PermutationsBasic_2_io_in_62_Im),
    .io_in_63_Re(PermutationsBasic_2_io_in_63_Re),
    .io_in_63_Im(PermutationsBasic_2_io_in_63_Im),
    .io_in_64_Re(PermutationsBasic_2_io_in_64_Re),
    .io_in_64_Im(PermutationsBasic_2_io_in_64_Im),
    .io_in_65_Re(PermutationsBasic_2_io_in_65_Re),
    .io_in_65_Im(PermutationsBasic_2_io_in_65_Im),
    .io_in_66_Re(PermutationsBasic_2_io_in_66_Re),
    .io_in_66_Im(PermutationsBasic_2_io_in_66_Im),
    .io_in_67_Re(PermutationsBasic_2_io_in_67_Re),
    .io_in_67_Im(PermutationsBasic_2_io_in_67_Im),
    .io_in_68_Re(PermutationsBasic_2_io_in_68_Re),
    .io_in_68_Im(PermutationsBasic_2_io_in_68_Im),
    .io_in_69_Re(PermutationsBasic_2_io_in_69_Re),
    .io_in_69_Im(PermutationsBasic_2_io_in_69_Im),
    .io_in_70_Re(PermutationsBasic_2_io_in_70_Re),
    .io_in_70_Im(PermutationsBasic_2_io_in_70_Im),
    .io_in_71_Re(PermutationsBasic_2_io_in_71_Re),
    .io_in_71_Im(PermutationsBasic_2_io_in_71_Im),
    .io_in_72_Re(PermutationsBasic_2_io_in_72_Re),
    .io_in_72_Im(PermutationsBasic_2_io_in_72_Im),
    .io_in_73_Re(PermutationsBasic_2_io_in_73_Re),
    .io_in_73_Im(PermutationsBasic_2_io_in_73_Im),
    .io_in_74_Re(PermutationsBasic_2_io_in_74_Re),
    .io_in_74_Im(PermutationsBasic_2_io_in_74_Im),
    .io_in_75_Re(PermutationsBasic_2_io_in_75_Re),
    .io_in_75_Im(PermutationsBasic_2_io_in_75_Im),
    .io_in_76_Re(PermutationsBasic_2_io_in_76_Re),
    .io_in_76_Im(PermutationsBasic_2_io_in_76_Im),
    .io_in_77_Re(PermutationsBasic_2_io_in_77_Re),
    .io_in_77_Im(PermutationsBasic_2_io_in_77_Im),
    .io_in_78_Re(PermutationsBasic_2_io_in_78_Re),
    .io_in_78_Im(PermutationsBasic_2_io_in_78_Im),
    .io_in_79_Re(PermutationsBasic_2_io_in_79_Re),
    .io_in_79_Im(PermutationsBasic_2_io_in_79_Im),
    .io_in_80_Re(PermutationsBasic_2_io_in_80_Re),
    .io_in_80_Im(PermutationsBasic_2_io_in_80_Im),
    .io_in_81_Re(PermutationsBasic_2_io_in_81_Re),
    .io_in_81_Im(PermutationsBasic_2_io_in_81_Im),
    .io_in_82_Re(PermutationsBasic_2_io_in_82_Re),
    .io_in_82_Im(PermutationsBasic_2_io_in_82_Im),
    .io_in_83_Re(PermutationsBasic_2_io_in_83_Re),
    .io_in_83_Im(PermutationsBasic_2_io_in_83_Im),
    .io_in_84_Re(PermutationsBasic_2_io_in_84_Re),
    .io_in_84_Im(PermutationsBasic_2_io_in_84_Im),
    .io_in_85_Re(PermutationsBasic_2_io_in_85_Re),
    .io_in_85_Im(PermutationsBasic_2_io_in_85_Im),
    .io_in_86_Re(PermutationsBasic_2_io_in_86_Re),
    .io_in_86_Im(PermutationsBasic_2_io_in_86_Im),
    .io_in_87_Re(PermutationsBasic_2_io_in_87_Re),
    .io_in_87_Im(PermutationsBasic_2_io_in_87_Im),
    .io_in_88_Re(PermutationsBasic_2_io_in_88_Re),
    .io_in_88_Im(PermutationsBasic_2_io_in_88_Im),
    .io_in_89_Re(PermutationsBasic_2_io_in_89_Re),
    .io_in_89_Im(PermutationsBasic_2_io_in_89_Im),
    .io_in_90_Re(PermutationsBasic_2_io_in_90_Re),
    .io_in_90_Im(PermutationsBasic_2_io_in_90_Im),
    .io_in_91_Re(PermutationsBasic_2_io_in_91_Re),
    .io_in_91_Im(PermutationsBasic_2_io_in_91_Im),
    .io_in_92_Re(PermutationsBasic_2_io_in_92_Re),
    .io_in_92_Im(PermutationsBasic_2_io_in_92_Im),
    .io_in_93_Re(PermutationsBasic_2_io_in_93_Re),
    .io_in_93_Im(PermutationsBasic_2_io_in_93_Im),
    .io_in_94_Re(PermutationsBasic_2_io_in_94_Re),
    .io_in_94_Im(PermutationsBasic_2_io_in_94_Im),
    .io_in_95_Re(PermutationsBasic_2_io_in_95_Re),
    .io_in_95_Im(PermutationsBasic_2_io_in_95_Im),
    .io_out_0_Re(PermutationsBasic_2_io_out_0_Re),
    .io_out_0_Im(PermutationsBasic_2_io_out_0_Im),
    .io_out_1_Re(PermutationsBasic_2_io_out_1_Re),
    .io_out_1_Im(PermutationsBasic_2_io_out_1_Im),
    .io_out_2_Re(PermutationsBasic_2_io_out_2_Re),
    .io_out_2_Im(PermutationsBasic_2_io_out_2_Im),
    .io_out_3_Re(PermutationsBasic_2_io_out_3_Re),
    .io_out_3_Im(PermutationsBasic_2_io_out_3_Im),
    .io_out_4_Re(PermutationsBasic_2_io_out_4_Re),
    .io_out_4_Im(PermutationsBasic_2_io_out_4_Im),
    .io_out_5_Re(PermutationsBasic_2_io_out_5_Re),
    .io_out_5_Im(PermutationsBasic_2_io_out_5_Im),
    .io_out_6_Re(PermutationsBasic_2_io_out_6_Re),
    .io_out_6_Im(PermutationsBasic_2_io_out_6_Im),
    .io_out_7_Re(PermutationsBasic_2_io_out_7_Re),
    .io_out_7_Im(PermutationsBasic_2_io_out_7_Im),
    .io_out_8_Re(PermutationsBasic_2_io_out_8_Re),
    .io_out_8_Im(PermutationsBasic_2_io_out_8_Im),
    .io_out_9_Re(PermutationsBasic_2_io_out_9_Re),
    .io_out_9_Im(PermutationsBasic_2_io_out_9_Im),
    .io_out_10_Re(PermutationsBasic_2_io_out_10_Re),
    .io_out_10_Im(PermutationsBasic_2_io_out_10_Im),
    .io_out_11_Re(PermutationsBasic_2_io_out_11_Re),
    .io_out_11_Im(PermutationsBasic_2_io_out_11_Im),
    .io_out_12_Re(PermutationsBasic_2_io_out_12_Re),
    .io_out_12_Im(PermutationsBasic_2_io_out_12_Im),
    .io_out_13_Re(PermutationsBasic_2_io_out_13_Re),
    .io_out_13_Im(PermutationsBasic_2_io_out_13_Im),
    .io_out_14_Re(PermutationsBasic_2_io_out_14_Re),
    .io_out_14_Im(PermutationsBasic_2_io_out_14_Im),
    .io_out_15_Re(PermutationsBasic_2_io_out_15_Re),
    .io_out_15_Im(PermutationsBasic_2_io_out_15_Im),
    .io_out_16_Re(PermutationsBasic_2_io_out_16_Re),
    .io_out_16_Im(PermutationsBasic_2_io_out_16_Im),
    .io_out_17_Re(PermutationsBasic_2_io_out_17_Re),
    .io_out_17_Im(PermutationsBasic_2_io_out_17_Im),
    .io_out_18_Re(PermutationsBasic_2_io_out_18_Re),
    .io_out_18_Im(PermutationsBasic_2_io_out_18_Im),
    .io_out_19_Re(PermutationsBasic_2_io_out_19_Re),
    .io_out_19_Im(PermutationsBasic_2_io_out_19_Im),
    .io_out_20_Re(PermutationsBasic_2_io_out_20_Re),
    .io_out_20_Im(PermutationsBasic_2_io_out_20_Im),
    .io_out_21_Re(PermutationsBasic_2_io_out_21_Re),
    .io_out_21_Im(PermutationsBasic_2_io_out_21_Im),
    .io_out_22_Re(PermutationsBasic_2_io_out_22_Re),
    .io_out_22_Im(PermutationsBasic_2_io_out_22_Im),
    .io_out_23_Re(PermutationsBasic_2_io_out_23_Re),
    .io_out_23_Im(PermutationsBasic_2_io_out_23_Im),
    .io_out_24_Re(PermutationsBasic_2_io_out_24_Re),
    .io_out_24_Im(PermutationsBasic_2_io_out_24_Im),
    .io_out_25_Re(PermutationsBasic_2_io_out_25_Re),
    .io_out_25_Im(PermutationsBasic_2_io_out_25_Im),
    .io_out_26_Re(PermutationsBasic_2_io_out_26_Re),
    .io_out_26_Im(PermutationsBasic_2_io_out_26_Im),
    .io_out_27_Re(PermutationsBasic_2_io_out_27_Re),
    .io_out_27_Im(PermutationsBasic_2_io_out_27_Im),
    .io_out_28_Re(PermutationsBasic_2_io_out_28_Re),
    .io_out_28_Im(PermutationsBasic_2_io_out_28_Im),
    .io_out_29_Re(PermutationsBasic_2_io_out_29_Re),
    .io_out_29_Im(PermutationsBasic_2_io_out_29_Im),
    .io_out_30_Re(PermutationsBasic_2_io_out_30_Re),
    .io_out_30_Im(PermutationsBasic_2_io_out_30_Im),
    .io_out_31_Re(PermutationsBasic_2_io_out_31_Re),
    .io_out_31_Im(PermutationsBasic_2_io_out_31_Im),
    .io_out_32_Re(PermutationsBasic_2_io_out_32_Re),
    .io_out_32_Im(PermutationsBasic_2_io_out_32_Im),
    .io_out_33_Re(PermutationsBasic_2_io_out_33_Re),
    .io_out_33_Im(PermutationsBasic_2_io_out_33_Im),
    .io_out_34_Re(PermutationsBasic_2_io_out_34_Re),
    .io_out_34_Im(PermutationsBasic_2_io_out_34_Im),
    .io_out_35_Re(PermutationsBasic_2_io_out_35_Re),
    .io_out_35_Im(PermutationsBasic_2_io_out_35_Im),
    .io_out_36_Re(PermutationsBasic_2_io_out_36_Re),
    .io_out_36_Im(PermutationsBasic_2_io_out_36_Im),
    .io_out_37_Re(PermutationsBasic_2_io_out_37_Re),
    .io_out_37_Im(PermutationsBasic_2_io_out_37_Im),
    .io_out_38_Re(PermutationsBasic_2_io_out_38_Re),
    .io_out_38_Im(PermutationsBasic_2_io_out_38_Im),
    .io_out_39_Re(PermutationsBasic_2_io_out_39_Re),
    .io_out_39_Im(PermutationsBasic_2_io_out_39_Im),
    .io_out_40_Re(PermutationsBasic_2_io_out_40_Re),
    .io_out_40_Im(PermutationsBasic_2_io_out_40_Im),
    .io_out_41_Re(PermutationsBasic_2_io_out_41_Re),
    .io_out_41_Im(PermutationsBasic_2_io_out_41_Im),
    .io_out_42_Re(PermutationsBasic_2_io_out_42_Re),
    .io_out_42_Im(PermutationsBasic_2_io_out_42_Im),
    .io_out_43_Re(PermutationsBasic_2_io_out_43_Re),
    .io_out_43_Im(PermutationsBasic_2_io_out_43_Im),
    .io_out_44_Re(PermutationsBasic_2_io_out_44_Re),
    .io_out_44_Im(PermutationsBasic_2_io_out_44_Im),
    .io_out_45_Re(PermutationsBasic_2_io_out_45_Re),
    .io_out_45_Im(PermutationsBasic_2_io_out_45_Im),
    .io_out_46_Re(PermutationsBasic_2_io_out_46_Re),
    .io_out_46_Im(PermutationsBasic_2_io_out_46_Im),
    .io_out_47_Re(PermutationsBasic_2_io_out_47_Re),
    .io_out_47_Im(PermutationsBasic_2_io_out_47_Im),
    .io_out_48_Re(PermutationsBasic_2_io_out_48_Re),
    .io_out_48_Im(PermutationsBasic_2_io_out_48_Im),
    .io_out_49_Re(PermutationsBasic_2_io_out_49_Re),
    .io_out_49_Im(PermutationsBasic_2_io_out_49_Im),
    .io_out_50_Re(PermutationsBasic_2_io_out_50_Re),
    .io_out_50_Im(PermutationsBasic_2_io_out_50_Im),
    .io_out_51_Re(PermutationsBasic_2_io_out_51_Re),
    .io_out_51_Im(PermutationsBasic_2_io_out_51_Im),
    .io_out_52_Re(PermutationsBasic_2_io_out_52_Re),
    .io_out_52_Im(PermutationsBasic_2_io_out_52_Im),
    .io_out_53_Re(PermutationsBasic_2_io_out_53_Re),
    .io_out_53_Im(PermutationsBasic_2_io_out_53_Im),
    .io_out_54_Re(PermutationsBasic_2_io_out_54_Re),
    .io_out_54_Im(PermutationsBasic_2_io_out_54_Im),
    .io_out_55_Re(PermutationsBasic_2_io_out_55_Re),
    .io_out_55_Im(PermutationsBasic_2_io_out_55_Im),
    .io_out_56_Re(PermutationsBasic_2_io_out_56_Re),
    .io_out_56_Im(PermutationsBasic_2_io_out_56_Im),
    .io_out_57_Re(PermutationsBasic_2_io_out_57_Re),
    .io_out_57_Im(PermutationsBasic_2_io_out_57_Im),
    .io_out_58_Re(PermutationsBasic_2_io_out_58_Re),
    .io_out_58_Im(PermutationsBasic_2_io_out_58_Im),
    .io_out_59_Re(PermutationsBasic_2_io_out_59_Re),
    .io_out_59_Im(PermutationsBasic_2_io_out_59_Im),
    .io_out_60_Re(PermutationsBasic_2_io_out_60_Re),
    .io_out_60_Im(PermutationsBasic_2_io_out_60_Im),
    .io_out_61_Re(PermutationsBasic_2_io_out_61_Re),
    .io_out_61_Im(PermutationsBasic_2_io_out_61_Im),
    .io_out_62_Re(PermutationsBasic_2_io_out_62_Re),
    .io_out_62_Im(PermutationsBasic_2_io_out_62_Im),
    .io_out_63_Re(PermutationsBasic_2_io_out_63_Re),
    .io_out_63_Im(PermutationsBasic_2_io_out_63_Im),
    .io_out_64_Re(PermutationsBasic_2_io_out_64_Re),
    .io_out_64_Im(PermutationsBasic_2_io_out_64_Im),
    .io_out_65_Re(PermutationsBasic_2_io_out_65_Re),
    .io_out_65_Im(PermutationsBasic_2_io_out_65_Im),
    .io_out_66_Re(PermutationsBasic_2_io_out_66_Re),
    .io_out_66_Im(PermutationsBasic_2_io_out_66_Im),
    .io_out_67_Re(PermutationsBasic_2_io_out_67_Re),
    .io_out_67_Im(PermutationsBasic_2_io_out_67_Im),
    .io_out_68_Re(PermutationsBasic_2_io_out_68_Re),
    .io_out_68_Im(PermutationsBasic_2_io_out_68_Im),
    .io_out_69_Re(PermutationsBasic_2_io_out_69_Re),
    .io_out_69_Im(PermutationsBasic_2_io_out_69_Im),
    .io_out_70_Re(PermutationsBasic_2_io_out_70_Re),
    .io_out_70_Im(PermutationsBasic_2_io_out_70_Im),
    .io_out_71_Re(PermutationsBasic_2_io_out_71_Re),
    .io_out_71_Im(PermutationsBasic_2_io_out_71_Im),
    .io_out_72_Re(PermutationsBasic_2_io_out_72_Re),
    .io_out_72_Im(PermutationsBasic_2_io_out_72_Im),
    .io_out_73_Re(PermutationsBasic_2_io_out_73_Re),
    .io_out_73_Im(PermutationsBasic_2_io_out_73_Im),
    .io_out_74_Re(PermutationsBasic_2_io_out_74_Re),
    .io_out_74_Im(PermutationsBasic_2_io_out_74_Im),
    .io_out_75_Re(PermutationsBasic_2_io_out_75_Re),
    .io_out_75_Im(PermutationsBasic_2_io_out_75_Im),
    .io_out_76_Re(PermutationsBasic_2_io_out_76_Re),
    .io_out_76_Im(PermutationsBasic_2_io_out_76_Im),
    .io_out_77_Re(PermutationsBasic_2_io_out_77_Re),
    .io_out_77_Im(PermutationsBasic_2_io_out_77_Im),
    .io_out_78_Re(PermutationsBasic_2_io_out_78_Re),
    .io_out_78_Im(PermutationsBasic_2_io_out_78_Im),
    .io_out_79_Re(PermutationsBasic_2_io_out_79_Re),
    .io_out_79_Im(PermutationsBasic_2_io_out_79_Im),
    .io_out_80_Re(PermutationsBasic_2_io_out_80_Re),
    .io_out_80_Im(PermutationsBasic_2_io_out_80_Im),
    .io_out_81_Re(PermutationsBasic_2_io_out_81_Re),
    .io_out_81_Im(PermutationsBasic_2_io_out_81_Im),
    .io_out_82_Re(PermutationsBasic_2_io_out_82_Re),
    .io_out_82_Im(PermutationsBasic_2_io_out_82_Im),
    .io_out_83_Re(PermutationsBasic_2_io_out_83_Re),
    .io_out_83_Im(PermutationsBasic_2_io_out_83_Im),
    .io_out_84_Re(PermutationsBasic_2_io_out_84_Re),
    .io_out_84_Im(PermutationsBasic_2_io_out_84_Im),
    .io_out_85_Re(PermutationsBasic_2_io_out_85_Re),
    .io_out_85_Im(PermutationsBasic_2_io_out_85_Im),
    .io_out_86_Re(PermutationsBasic_2_io_out_86_Re),
    .io_out_86_Im(PermutationsBasic_2_io_out_86_Im),
    .io_out_87_Re(PermutationsBasic_2_io_out_87_Re),
    .io_out_87_Im(PermutationsBasic_2_io_out_87_Im),
    .io_out_88_Re(PermutationsBasic_2_io_out_88_Re),
    .io_out_88_Im(PermutationsBasic_2_io_out_88_Im),
    .io_out_89_Re(PermutationsBasic_2_io_out_89_Re),
    .io_out_89_Im(PermutationsBasic_2_io_out_89_Im),
    .io_out_90_Re(PermutationsBasic_2_io_out_90_Re),
    .io_out_90_Im(PermutationsBasic_2_io_out_90_Im),
    .io_out_91_Re(PermutationsBasic_2_io_out_91_Re),
    .io_out_91_Im(PermutationsBasic_2_io_out_91_Im),
    .io_out_92_Re(PermutationsBasic_2_io_out_92_Re),
    .io_out_92_Im(PermutationsBasic_2_io_out_92_Im),
    .io_out_93_Re(PermutationsBasic_2_io_out_93_Re),
    .io_out_93_Im(PermutationsBasic_2_io_out_93_Im),
    .io_out_94_Re(PermutationsBasic_2_io_out_94_Re),
    .io_out_94_Im(PermutationsBasic_2_io_out_94_Im),
    .io_out_95_Re(PermutationsBasic_2_io_out_95_Re),
    .io_out_95_Im(PermutationsBasic_2_io_out_95_Im)
  );
  TwiddleFactors_mr TwiddleFactors_mr ( // @[FFTDesigns.scala 3454:29]
    .clock(TwiddleFactors_mr_clock),
    .reset(TwiddleFactors_mr_reset),
    .io_in_0_Re(TwiddleFactors_mr_io_in_0_Re),
    .io_in_0_Im(TwiddleFactors_mr_io_in_0_Im),
    .io_in_1_Re(TwiddleFactors_mr_io_in_1_Re),
    .io_in_1_Im(TwiddleFactors_mr_io_in_1_Im),
    .io_in_2_Re(TwiddleFactors_mr_io_in_2_Re),
    .io_in_2_Im(TwiddleFactors_mr_io_in_2_Im),
    .io_in_3_Re(TwiddleFactors_mr_io_in_3_Re),
    .io_in_3_Im(TwiddleFactors_mr_io_in_3_Im),
    .io_in_4_Re(TwiddleFactors_mr_io_in_4_Re),
    .io_in_4_Im(TwiddleFactors_mr_io_in_4_Im),
    .io_in_5_Re(TwiddleFactors_mr_io_in_5_Re),
    .io_in_5_Im(TwiddleFactors_mr_io_in_5_Im),
    .io_in_6_Re(TwiddleFactors_mr_io_in_6_Re),
    .io_in_6_Im(TwiddleFactors_mr_io_in_6_Im),
    .io_in_7_Re(TwiddleFactors_mr_io_in_7_Re),
    .io_in_7_Im(TwiddleFactors_mr_io_in_7_Im),
    .io_in_8_Re(TwiddleFactors_mr_io_in_8_Re),
    .io_in_8_Im(TwiddleFactors_mr_io_in_8_Im),
    .io_in_9_Re(TwiddleFactors_mr_io_in_9_Re),
    .io_in_9_Im(TwiddleFactors_mr_io_in_9_Im),
    .io_in_10_Re(TwiddleFactors_mr_io_in_10_Re),
    .io_in_10_Im(TwiddleFactors_mr_io_in_10_Im),
    .io_in_11_Re(TwiddleFactors_mr_io_in_11_Re),
    .io_in_11_Im(TwiddleFactors_mr_io_in_11_Im),
    .io_in_12_Re(TwiddleFactors_mr_io_in_12_Re),
    .io_in_12_Im(TwiddleFactors_mr_io_in_12_Im),
    .io_in_13_Re(TwiddleFactors_mr_io_in_13_Re),
    .io_in_13_Im(TwiddleFactors_mr_io_in_13_Im),
    .io_in_14_Re(TwiddleFactors_mr_io_in_14_Re),
    .io_in_14_Im(TwiddleFactors_mr_io_in_14_Im),
    .io_in_15_Re(TwiddleFactors_mr_io_in_15_Re),
    .io_in_15_Im(TwiddleFactors_mr_io_in_15_Im),
    .io_in_16_Re(TwiddleFactors_mr_io_in_16_Re),
    .io_in_16_Im(TwiddleFactors_mr_io_in_16_Im),
    .io_in_17_Re(TwiddleFactors_mr_io_in_17_Re),
    .io_in_17_Im(TwiddleFactors_mr_io_in_17_Im),
    .io_in_18_Re(TwiddleFactors_mr_io_in_18_Re),
    .io_in_18_Im(TwiddleFactors_mr_io_in_18_Im),
    .io_in_19_Re(TwiddleFactors_mr_io_in_19_Re),
    .io_in_19_Im(TwiddleFactors_mr_io_in_19_Im),
    .io_in_20_Re(TwiddleFactors_mr_io_in_20_Re),
    .io_in_20_Im(TwiddleFactors_mr_io_in_20_Im),
    .io_in_21_Re(TwiddleFactors_mr_io_in_21_Re),
    .io_in_21_Im(TwiddleFactors_mr_io_in_21_Im),
    .io_in_22_Re(TwiddleFactors_mr_io_in_22_Re),
    .io_in_22_Im(TwiddleFactors_mr_io_in_22_Im),
    .io_in_23_Re(TwiddleFactors_mr_io_in_23_Re),
    .io_in_23_Im(TwiddleFactors_mr_io_in_23_Im),
    .io_in_24_Re(TwiddleFactors_mr_io_in_24_Re),
    .io_in_24_Im(TwiddleFactors_mr_io_in_24_Im),
    .io_in_25_Re(TwiddleFactors_mr_io_in_25_Re),
    .io_in_25_Im(TwiddleFactors_mr_io_in_25_Im),
    .io_in_26_Re(TwiddleFactors_mr_io_in_26_Re),
    .io_in_26_Im(TwiddleFactors_mr_io_in_26_Im),
    .io_in_27_Re(TwiddleFactors_mr_io_in_27_Re),
    .io_in_27_Im(TwiddleFactors_mr_io_in_27_Im),
    .io_in_28_Re(TwiddleFactors_mr_io_in_28_Re),
    .io_in_28_Im(TwiddleFactors_mr_io_in_28_Im),
    .io_in_29_Re(TwiddleFactors_mr_io_in_29_Re),
    .io_in_29_Im(TwiddleFactors_mr_io_in_29_Im),
    .io_in_30_Re(TwiddleFactors_mr_io_in_30_Re),
    .io_in_30_Im(TwiddleFactors_mr_io_in_30_Im),
    .io_in_31_Re(TwiddleFactors_mr_io_in_31_Re),
    .io_in_31_Im(TwiddleFactors_mr_io_in_31_Im),
    .io_in_32_Re(TwiddleFactors_mr_io_in_32_Re),
    .io_in_32_Im(TwiddleFactors_mr_io_in_32_Im),
    .io_in_33_Re(TwiddleFactors_mr_io_in_33_Re),
    .io_in_33_Im(TwiddleFactors_mr_io_in_33_Im),
    .io_in_34_Re(TwiddleFactors_mr_io_in_34_Re),
    .io_in_34_Im(TwiddleFactors_mr_io_in_34_Im),
    .io_in_35_Re(TwiddleFactors_mr_io_in_35_Re),
    .io_in_35_Im(TwiddleFactors_mr_io_in_35_Im),
    .io_in_36_Re(TwiddleFactors_mr_io_in_36_Re),
    .io_in_36_Im(TwiddleFactors_mr_io_in_36_Im),
    .io_in_37_Re(TwiddleFactors_mr_io_in_37_Re),
    .io_in_37_Im(TwiddleFactors_mr_io_in_37_Im),
    .io_in_38_Re(TwiddleFactors_mr_io_in_38_Re),
    .io_in_38_Im(TwiddleFactors_mr_io_in_38_Im),
    .io_in_39_Re(TwiddleFactors_mr_io_in_39_Re),
    .io_in_39_Im(TwiddleFactors_mr_io_in_39_Im),
    .io_in_40_Re(TwiddleFactors_mr_io_in_40_Re),
    .io_in_40_Im(TwiddleFactors_mr_io_in_40_Im),
    .io_in_41_Re(TwiddleFactors_mr_io_in_41_Re),
    .io_in_41_Im(TwiddleFactors_mr_io_in_41_Im),
    .io_in_42_Re(TwiddleFactors_mr_io_in_42_Re),
    .io_in_42_Im(TwiddleFactors_mr_io_in_42_Im),
    .io_in_43_Re(TwiddleFactors_mr_io_in_43_Re),
    .io_in_43_Im(TwiddleFactors_mr_io_in_43_Im),
    .io_in_44_Re(TwiddleFactors_mr_io_in_44_Re),
    .io_in_44_Im(TwiddleFactors_mr_io_in_44_Im),
    .io_in_45_Re(TwiddleFactors_mr_io_in_45_Re),
    .io_in_45_Im(TwiddleFactors_mr_io_in_45_Im),
    .io_in_46_Re(TwiddleFactors_mr_io_in_46_Re),
    .io_in_46_Im(TwiddleFactors_mr_io_in_46_Im),
    .io_in_47_Re(TwiddleFactors_mr_io_in_47_Re),
    .io_in_47_Im(TwiddleFactors_mr_io_in_47_Im),
    .io_in_48_Re(TwiddleFactors_mr_io_in_48_Re),
    .io_in_48_Im(TwiddleFactors_mr_io_in_48_Im),
    .io_in_49_Re(TwiddleFactors_mr_io_in_49_Re),
    .io_in_49_Im(TwiddleFactors_mr_io_in_49_Im),
    .io_in_50_Re(TwiddleFactors_mr_io_in_50_Re),
    .io_in_50_Im(TwiddleFactors_mr_io_in_50_Im),
    .io_in_51_Re(TwiddleFactors_mr_io_in_51_Re),
    .io_in_51_Im(TwiddleFactors_mr_io_in_51_Im),
    .io_in_52_Re(TwiddleFactors_mr_io_in_52_Re),
    .io_in_52_Im(TwiddleFactors_mr_io_in_52_Im),
    .io_in_53_Re(TwiddleFactors_mr_io_in_53_Re),
    .io_in_53_Im(TwiddleFactors_mr_io_in_53_Im),
    .io_in_54_Re(TwiddleFactors_mr_io_in_54_Re),
    .io_in_54_Im(TwiddleFactors_mr_io_in_54_Im),
    .io_in_55_Re(TwiddleFactors_mr_io_in_55_Re),
    .io_in_55_Im(TwiddleFactors_mr_io_in_55_Im),
    .io_in_56_Re(TwiddleFactors_mr_io_in_56_Re),
    .io_in_56_Im(TwiddleFactors_mr_io_in_56_Im),
    .io_in_57_Re(TwiddleFactors_mr_io_in_57_Re),
    .io_in_57_Im(TwiddleFactors_mr_io_in_57_Im),
    .io_in_58_Re(TwiddleFactors_mr_io_in_58_Re),
    .io_in_58_Im(TwiddleFactors_mr_io_in_58_Im),
    .io_in_59_Re(TwiddleFactors_mr_io_in_59_Re),
    .io_in_59_Im(TwiddleFactors_mr_io_in_59_Im),
    .io_in_60_Re(TwiddleFactors_mr_io_in_60_Re),
    .io_in_60_Im(TwiddleFactors_mr_io_in_60_Im),
    .io_in_61_Re(TwiddleFactors_mr_io_in_61_Re),
    .io_in_61_Im(TwiddleFactors_mr_io_in_61_Im),
    .io_in_62_Re(TwiddleFactors_mr_io_in_62_Re),
    .io_in_62_Im(TwiddleFactors_mr_io_in_62_Im),
    .io_in_63_Re(TwiddleFactors_mr_io_in_63_Re),
    .io_in_63_Im(TwiddleFactors_mr_io_in_63_Im),
    .io_in_64_Re(TwiddleFactors_mr_io_in_64_Re),
    .io_in_64_Im(TwiddleFactors_mr_io_in_64_Im),
    .io_in_65_Re(TwiddleFactors_mr_io_in_65_Re),
    .io_in_65_Im(TwiddleFactors_mr_io_in_65_Im),
    .io_in_66_Re(TwiddleFactors_mr_io_in_66_Re),
    .io_in_66_Im(TwiddleFactors_mr_io_in_66_Im),
    .io_in_67_Re(TwiddleFactors_mr_io_in_67_Re),
    .io_in_67_Im(TwiddleFactors_mr_io_in_67_Im),
    .io_in_68_Re(TwiddleFactors_mr_io_in_68_Re),
    .io_in_68_Im(TwiddleFactors_mr_io_in_68_Im),
    .io_in_69_Re(TwiddleFactors_mr_io_in_69_Re),
    .io_in_69_Im(TwiddleFactors_mr_io_in_69_Im),
    .io_in_70_Re(TwiddleFactors_mr_io_in_70_Re),
    .io_in_70_Im(TwiddleFactors_mr_io_in_70_Im),
    .io_in_71_Re(TwiddleFactors_mr_io_in_71_Re),
    .io_in_71_Im(TwiddleFactors_mr_io_in_71_Im),
    .io_in_72_Re(TwiddleFactors_mr_io_in_72_Re),
    .io_in_72_Im(TwiddleFactors_mr_io_in_72_Im),
    .io_in_73_Re(TwiddleFactors_mr_io_in_73_Re),
    .io_in_73_Im(TwiddleFactors_mr_io_in_73_Im),
    .io_in_74_Re(TwiddleFactors_mr_io_in_74_Re),
    .io_in_74_Im(TwiddleFactors_mr_io_in_74_Im),
    .io_in_75_Re(TwiddleFactors_mr_io_in_75_Re),
    .io_in_75_Im(TwiddleFactors_mr_io_in_75_Im),
    .io_in_76_Re(TwiddleFactors_mr_io_in_76_Re),
    .io_in_76_Im(TwiddleFactors_mr_io_in_76_Im),
    .io_in_77_Re(TwiddleFactors_mr_io_in_77_Re),
    .io_in_77_Im(TwiddleFactors_mr_io_in_77_Im),
    .io_in_78_Re(TwiddleFactors_mr_io_in_78_Re),
    .io_in_78_Im(TwiddleFactors_mr_io_in_78_Im),
    .io_in_79_Re(TwiddleFactors_mr_io_in_79_Re),
    .io_in_79_Im(TwiddleFactors_mr_io_in_79_Im),
    .io_in_80_Re(TwiddleFactors_mr_io_in_80_Re),
    .io_in_80_Im(TwiddleFactors_mr_io_in_80_Im),
    .io_in_81_Re(TwiddleFactors_mr_io_in_81_Re),
    .io_in_81_Im(TwiddleFactors_mr_io_in_81_Im),
    .io_in_82_Re(TwiddleFactors_mr_io_in_82_Re),
    .io_in_82_Im(TwiddleFactors_mr_io_in_82_Im),
    .io_in_83_Re(TwiddleFactors_mr_io_in_83_Re),
    .io_in_83_Im(TwiddleFactors_mr_io_in_83_Im),
    .io_in_84_Re(TwiddleFactors_mr_io_in_84_Re),
    .io_in_84_Im(TwiddleFactors_mr_io_in_84_Im),
    .io_in_85_Re(TwiddleFactors_mr_io_in_85_Re),
    .io_in_85_Im(TwiddleFactors_mr_io_in_85_Im),
    .io_in_86_Re(TwiddleFactors_mr_io_in_86_Re),
    .io_in_86_Im(TwiddleFactors_mr_io_in_86_Im),
    .io_in_87_Re(TwiddleFactors_mr_io_in_87_Re),
    .io_in_87_Im(TwiddleFactors_mr_io_in_87_Im),
    .io_in_88_Re(TwiddleFactors_mr_io_in_88_Re),
    .io_in_88_Im(TwiddleFactors_mr_io_in_88_Im),
    .io_in_89_Re(TwiddleFactors_mr_io_in_89_Re),
    .io_in_89_Im(TwiddleFactors_mr_io_in_89_Im),
    .io_in_90_Re(TwiddleFactors_mr_io_in_90_Re),
    .io_in_90_Im(TwiddleFactors_mr_io_in_90_Im),
    .io_in_91_Re(TwiddleFactors_mr_io_in_91_Re),
    .io_in_91_Im(TwiddleFactors_mr_io_in_91_Im),
    .io_in_92_Re(TwiddleFactors_mr_io_in_92_Re),
    .io_in_92_Im(TwiddleFactors_mr_io_in_92_Im),
    .io_in_93_Re(TwiddleFactors_mr_io_in_93_Re),
    .io_in_93_Im(TwiddleFactors_mr_io_in_93_Im),
    .io_in_94_Re(TwiddleFactors_mr_io_in_94_Re),
    .io_in_94_Im(TwiddleFactors_mr_io_in_94_Im),
    .io_in_95_Re(TwiddleFactors_mr_io_in_95_Re),
    .io_in_95_Im(TwiddleFactors_mr_io_in_95_Im),
    .io_out_0_Re(TwiddleFactors_mr_io_out_0_Re),
    .io_out_0_Im(TwiddleFactors_mr_io_out_0_Im),
    .io_out_1_Re(TwiddleFactors_mr_io_out_1_Re),
    .io_out_1_Im(TwiddleFactors_mr_io_out_1_Im),
    .io_out_2_Re(TwiddleFactors_mr_io_out_2_Re),
    .io_out_2_Im(TwiddleFactors_mr_io_out_2_Im),
    .io_out_3_Re(TwiddleFactors_mr_io_out_3_Re),
    .io_out_3_Im(TwiddleFactors_mr_io_out_3_Im),
    .io_out_4_Re(TwiddleFactors_mr_io_out_4_Re),
    .io_out_4_Im(TwiddleFactors_mr_io_out_4_Im),
    .io_out_5_Re(TwiddleFactors_mr_io_out_5_Re),
    .io_out_5_Im(TwiddleFactors_mr_io_out_5_Im),
    .io_out_6_Re(TwiddleFactors_mr_io_out_6_Re),
    .io_out_6_Im(TwiddleFactors_mr_io_out_6_Im),
    .io_out_7_Re(TwiddleFactors_mr_io_out_7_Re),
    .io_out_7_Im(TwiddleFactors_mr_io_out_7_Im),
    .io_out_8_Re(TwiddleFactors_mr_io_out_8_Re),
    .io_out_8_Im(TwiddleFactors_mr_io_out_8_Im),
    .io_out_9_Re(TwiddleFactors_mr_io_out_9_Re),
    .io_out_9_Im(TwiddleFactors_mr_io_out_9_Im),
    .io_out_10_Re(TwiddleFactors_mr_io_out_10_Re),
    .io_out_10_Im(TwiddleFactors_mr_io_out_10_Im),
    .io_out_11_Re(TwiddleFactors_mr_io_out_11_Re),
    .io_out_11_Im(TwiddleFactors_mr_io_out_11_Im),
    .io_out_12_Re(TwiddleFactors_mr_io_out_12_Re),
    .io_out_12_Im(TwiddleFactors_mr_io_out_12_Im),
    .io_out_13_Re(TwiddleFactors_mr_io_out_13_Re),
    .io_out_13_Im(TwiddleFactors_mr_io_out_13_Im),
    .io_out_14_Re(TwiddleFactors_mr_io_out_14_Re),
    .io_out_14_Im(TwiddleFactors_mr_io_out_14_Im),
    .io_out_15_Re(TwiddleFactors_mr_io_out_15_Re),
    .io_out_15_Im(TwiddleFactors_mr_io_out_15_Im),
    .io_out_16_Re(TwiddleFactors_mr_io_out_16_Re),
    .io_out_16_Im(TwiddleFactors_mr_io_out_16_Im),
    .io_out_17_Re(TwiddleFactors_mr_io_out_17_Re),
    .io_out_17_Im(TwiddleFactors_mr_io_out_17_Im),
    .io_out_18_Re(TwiddleFactors_mr_io_out_18_Re),
    .io_out_18_Im(TwiddleFactors_mr_io_out_18_Im),
    .io_out_19_Re(TwiddleFactors_mr_io_out_19_Re),
    .io_out_19_Im(TwiddleFactors_mr_io_out_19_Im),
    .io_out_20_Re(TwiddleFactors_mr_io_out_20_Re),
    .io_out_20_Im(TwiddleFactors_mr_io_out_20_Im),
    .io_out_21_Re(TwiddleFactors_mr_io_out_21_Re),
    .io_out_21_Im(TwiddleFactors_mr_io_out_21_Im),
    .io_out_22_Re(TwiddleFactors_mr_io_out_22_Re),
    .io_out_22_Im(TwiddleFactors_mr_io_out_22_Im),
    .io_out_23_Re(TwiddleFactors_mr_io_out_23_Re),
    .io_out_23_Im(TwiddleFactors_mr_io_out_23_Im),
    .io_out_24_Re(TwiddleFactors_mr_io_out_24_Re),
    .io_out_24_Im(TwiddleFactors_mr_io_out_24_Im),
    .io_out_25_Re(TwiddleFactors_mr_io_out_25_Re),
    .io_out_25_Im(TwiddleFactors_mr_io_out_25_Im),
    .io_out_26_Re(TwiddleFactors_mr_io_out_26_Re),
    .io_out_26_Im(TwiddleFactors_mr_io_out_26_Im),
    .io_out_27_Re(TwiddleFactors_mr_io_out_27_Re),
    .io_out_27_Im(TwiddleFactors_mr_io_out_27_Im),
    .io_out_28_Re(TwiddleFactors_mr_io_out_28_Re),
    .io_out_28_Im(TwiddleFactors_mr_io_out_28_Im),
    .io_out_29_Re(TwiddleFactors_mr_io_out_29_Re),
    .io_out_29_Im(TwiddleFactors_mr_io_out_29_Im),
    .io_out_30_Re(TwiddleFactors_mr_io_out_30_Re),
    .io_out_30_Im(TwiddleFactors_mr_io_out_30_Im),
    .io_out_31_Re(TwiddleFactors_mr_io_out_31_Re),
    .io_out_31_Im(TwiddleFactors_mr_io_out_31_Im),
    .io_out_32_Re(TwiddleFactors_mr_io_out_32_Re),
    .io_out_32_Im(TwiddleFactors_mr_io_out_32_Im),
    .io_out_33_Re(TwiddleFactors_mr_io_out_33_Re),
    .io_out_33_Im(TwiddleFactors_mr_io_out_33_Im),
    .io_out_34_Re(TwiddleFactors_mr_io_out_34_Re),
    .io_out_34_Im(TwiddleFactors_mr_io_out_34_Im),
    .io_out_35_Re(TwiddleFactors_mr_io_out_35_Re),
    .io_out_35_Im(TwiddleFactors_mr_io_out_35_Im),
    .io_out_36_Re(TwiddleFactors_mr_io_out_36_Re),
    .io_out_36_Im(TwiddleFactors_mr_io_out_36_Im),
    .io_out_37_Re(TwiddleFactors_mr_io_out_37_Re),
    .io_out_37_Im(TwiddleFactors_mr_io_out_37_Im),
    .io_out_38_Re(TwiddleFactors_mr_io_out_38_Re),
    .io_out_38_Im(TwiddleFactors_mr_io_out_38_Im),
    .io_out_39_Re(TwiddleFactors_mr_io_out_39_Re),
    .io_out_39_Im(TwiddleFactors_mr_io_out_39_Im),
    .io_out_40_Re(TwiddleFactors_mr_io_out_40_Re),
    .io_out_40_Im(TwiddleFactors_mr_io_out_40_Im),
    .io_out_41_Re(TwiddleFactors_mr_io_out_41_Re),
    .io_out_41_Im(TwiddleFactors_mr_io_out_41_Im),
    .io_out_42_Re(TwiddleFactors_mr_io_out_42_Re),
    .io_out_42_Im(TwiddleFactors_mr_io_out_42_Im),
    .io_out_43_Re(TwiddleFactors_mr_io_out_43_Re),
    .io_out_43_Im(TwiddleFactors_mr_io_out_43_Im),
    .io_out_44_Re(TwiddleFactors_mr_io_out_44_Re),
    .io_out_44_Im(TwiddleFactors_mr_io_out_44_Im),
    .io_out_45_Re(TwiddleFactors_mr_io_out_45_Re),
    .io_out_45_Im(TwiddleFactors_mr_io_out_45_Im),
    .io_out_46_Re(TwiddleFactors_mr_io_out_46_Re),
    .io_out_46_Im(TwiddleFactors_mr_io_out_46_Im),
    .io_out_47_Re(TwiddleFactors_mr_io_out_47_Re),
    .io_out_47_Im(TwiddleFactors_mr_io_out_47_Im),
    .io_out_48_Re(TwiddleFactors_mr_io_out_48_Re),
    .io_out_48_Im(TwiddleFactors_mr_io_out_48_Im),
    .io_out_49_Re(TwiddleFactors_mr_io_out_49_Re),
    .io_out_49_Im(TwiddleFactors_mr_io_out_49_Im),
    .io_out_50_Re(TwiddleFactors_mr_io_out_50_Re),
    .io_out_50_Im(TwiddleFactors_mr_io_out_50_Im),
    .io_out_51_Re(TwiddleFactors_mr_io_out_51_Re),
    .io_out_51_Im(TwiddleFactors_mr_io_out_51_Im),
    .io_out_52_Re(TwiddleFactors_mr_io_out_52_Re),
    .io_out_52_Im(TwiddleFactors_mr_io_out_52_Im),
    .io_out_53_Re(TwiddleFactors_mr_io_out_53_Re),
    .io_out_53_Im(TwiddleFactors_mr_io_out_53_Im),
    .io_out_54_Re(TwiddleFactors_mr_io_out_54_Re),
    .io_out_54_Im(TwiddleFactors_mr_io_out_54_Im),
    .io_out_55_Re(TwiddleFactors_mr_io_out_55_Re),
    .io_out_55_Im(TwiddleFactors_mr_io_out_55_Im),
    .io_out_56_Re(TwiddleFactors_mr_io_out_56_Re),
    .io_out_56_Im(TwiddleFactors_mr_io_out_56_Im),
    .io_out_57_Re(TwiddleFactors_mr_io_out_57_Re),
    .io_out_57_Im(TwiddleFactors_mr_io_out_57_Im),
    .io_out_58_Re(TwiddleFactors_mr_io_out_58_Re),
    .io_out_58_Im(TwiddleFactors_mr_io_out_58_Im),
    .io_out_59_Re(TwiddleFactors_mr_io_out_59_Re),
    .io_out_59_Im(TwiddleFactors_mr_io_out_59_Im),
    .io_out_60_Re(TwiddleFactors_mr_io_out_60_Re),
    .io_out_60_Im(TwiddleFactors_mr_io_out_60_Im),
    .io_out_61_Re(TwiddleFactors_mr_io_out_61_Re),
    .io_out_61_Im(TwiddleFactors_mr_io_out_61_Im),
    .io_out_62_Re(TwiddleFactors_mr_io_out_62_Re),
    .io_out_62_Im(TwiddleFactors_mr_io_out_62_Im),
    .io_out_63_Re(TwiddleFactors_mr_io_out_63_Re),
    .io_out_63_Im(TwiddleFactors_mr_io_out_63_Im),
    .io_out_64_Re(TwiddleFactors_mr_io_out_64_Re),
    .io_out_64_Im(TwiddleFactors_mr_io_out_64_Im),
    .io_out_65_Re(TwiddleFactors_mr_io_out_65_Re),
    .io_out_65_Im(TwiddleFactors_mr_io_out_65_Im),
    .io_out_66_Re(TwiddleFactors_mr_io_out_66_Re),
    .io_out_66_Im(TwiddleFactors_mr_io_out_66_Im),
    .io_out_67_Re(TwiddleFactors_mr_io_out_67_Re),
    .io_out_67_Im(TwiddleFactors_mr_io_out_67_Im),
    .io_out_68_Re(TwiddleFactors_mr_io_out_68_Re),
    .io_out_68_Im(TwiddleFactors_mr_io_out_68_Im),
    .io_out_69_Re(TwiddleFactors_mr_io_out_69_Re),
    .io_out_69_Im(TwiddleFactors_mr_io_out_69_Im),
    .io_out_70_Re(TwiddleFactors_mr_io_out_70_Re),
    .io_out_70_Im(TwiddleFactors_mr_io_out_70_Im),
    .io_out_71_Re(TwiddleFactors_mr_io_out_71_Re),
    .io_out_71_Im(TwiddleFactors_mr_io_out_71_Im),
    .io_out_72_Re(TwiddleFactors_mr_io_out_72_Re),
    .io_out_72_Im(TwiddleFactors_mr_io_out_72_Im),
    .io_out_73_Re(TwiddleFactors_mr_io_out_73_Re),
    .io_out_73_Im(TwiddleFactors_mr_io_out_73_Im),
    .io_out_74_Re(TwiddleFactors_mr_io_out_74_Re),
    .io_out_74_Im(TwiddleFactors_mr_io_out_74_Im),
    .io_out_75_Re(TwiddleFactors_mr_io_out_75_Re),
    .io_out_75_Im(TwiddleFactors_mr_io_out_75_Im),
    .io_out_76_Re(TwiddleFactors_mr_io_out_76_Re),
    .io_out_76_Im(TwiddleFactors_mr_io_out_76_Im),
    .io_out_77_Re(TwiddleFactors_mr_io_out_77_Re),
    .io_out_77_Im(TwiddleFactors_mr_io_out_77_Im),
    .io_out_78_Re(TwiddleFactors_mr_io_out_78_Re),
    .io_out_78_Im(TwiddleFactors_mr_io_out_78_Im),
    .io_out_79_Re(TwiddleFactors_mr_io_out_79_Re),
    .io_out_79_Im(TwiddleFactors_mr_io_out_79_Im),
    .io_out_80_Re(TwiddleFactors_mr_io_out_80_Re),
    .io_out_80_Im(TwiddleFactors_mr_io_out_80_Im),
    .io_out_81_Re(TwiddleFactors_mr_io_out_81_Re),
    .io_out_81_Im(TwiddleFactors_mr_io_out_81_Im),
    .io_out_82_Re(TwiddleFactors_mr_io_out_82_Re),
    .io_out_82_Im(TwiddleFactors_mr_io_out_82_Im),
    .io_out_83_Re(TwiddleFactors_mr_io_out_83_Re),
    .io_out_83_Im(TwiddleFactors_mr_io_out_83_Im),
    .io_out_84_Re(TwiddleFactors_mr_io_out_84_Re),
    .io_out_84_Im(TwiddleFactors_mr_io_out_84_Im),
    .io_out_85_Re(TwiddleFactors_mr_io_out_85_Re),
    .io_out_85_Im(TwiddleFactors_mr_io_out_85_Im),
    .io_out_86_Re(TwiddleFactors_mr_io_out_86_Re),
    .io_out_86_Im(TwiddleFactors_mr_io_out_86_Im),
    .io_out_87_Re(TwiddleFactors_mr_io_out_87_Re),
    .io_out_87_Im(TwiddleFactors_mr_io_out_87_Im),
    .io_out_88_Re(TwiddleFactors_mr_io_out_88_Re),
    .io_out_88_Im(TwiddleFactors_mr_io_out_88_Im),
    .io_out_89_Re(TwiddleFactors_mr_io_out_89_Re),
    .io_out_89_Im(TwiddleFactors_mr_io_out_89_Im),
    .io_out_90_Re(TwiddleFactors_mr_io_out_90_Re),
    .io_out_90_Im(TwiddleFactors_mr_io_out_90_Im),
    .io_out_91_Re(TwiddleFactors_mr_io_out_91_Re),
    .io_out_91_Im(TwiddleFactors_mr_io_out_91_Im),
    .io_out_92_Re(TwiddleFactors_mr_io_out_92_Re),
    .io_out_92_Im(TwiddleFactors_mr_io_out_92_Im),
    .io_out_93_Re(TwiddleFactors_mr_io_out_93_Re),
    .io_out_93_Im(TwiddleFactors_mr_io_out_93_Im),
    .io_out_94_Re(TwiddleFactors_mr_io_out_94_Re),
    .io_out_94_Im(TwiddleFactors_mr_io_out_94_Im),
    .io_out_95_Re(TwiddleFactors_mr_io_out_95_Re),
    .io_out_95_Im(TwiddleFactors_mr_io_out_95_Im)
  );
  assign io_out_validate = out_regdelay; // @[FFTDesigns.scala 3473:21]
  assign io_out_0_Re = out_results_0_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_0_Im = out_results_0_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_1_Re = out_results_1_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_1_Im = out_results_1_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_2_Re = out_results_2_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_2_Im = out_results_2_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_3_Re = out_results_3_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_3_Im = out_results_3_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_4_Re = out_results_4_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_4_Im = out_results_4_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_5_Re = out_results_5_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_5_Im = out_results_5_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_6_Re = out_results_6_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_6_Im = out_results_6_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_7_Re = out_results_7_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_7_Im = out_results_7_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_8_Re = out_results_8_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_8_Im = out_results_8_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_9_Re = out_results_9_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_9_Im = out_results_9_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_10_Re = out_results_10_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_10_Im = out_results_10_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_11_Re = out_results_11_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_11_Im = out_results_11_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_12_Re = out_results_12_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_12_Im = out_results_12_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_13_Re = out_results_13_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_13_Im = out_results_13_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_14_Re = out_results_14_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_14_Im = out_results_14_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_15_Re = out_results_15_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_15_Im = out_results_15_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_16_Re = out_results_16_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_16_Im = out_results_16_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_17_Re = out_results_17_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_17_Im = out_results_17_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_18_Re = out_results_18_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_18_Im = out_results_18_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_19_Re = out_results_19_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_19_Im = out_results_19_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_20_Re = out_results_20_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_20_Im = out_results_20_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_21_Re = out_results_21_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_21_Im = out_results_21_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_22_Re = out_results_22_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_22_Im = out_results_22_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_23_Re = out_results_23_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_23_Im = out_results_23_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_24_Re = out_results_24_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_24_Im = out_results_24_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_25_Re = out_results_25_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_25_Im = out_results_25_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_26_Re = out_results_26_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_26_Im = out_results_26_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_27_Re = out_results_27_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_27_Im = out_results_27_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_28_Re = out_results_28_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_28_Im = out_results_28_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_29_Re = out_results_29_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_29_Im = out_results_29_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_30_Re = out_results_30_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_30_Im = out_results_30_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_31_Re = out_results_31_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_31_Im = out_results_31_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_32_Re = out_results_32_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_32_Im = out_results_32_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_33_Re = out_results_33_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_33_Im = out_results_33_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_34_Re = out_results_34_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_34_Im = out_results_34_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_35_Re = out_results_35_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_35_Im = out_results_35_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_36_Re = out_results_36_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_36_Im = out_results_36_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_37_Re = out_results_37_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_37_Im = out_results_37_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_38_Re = out_results_38_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_38_Im = out_results_38_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_39_Re = out_results_39_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_39_Im = out_results_39_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_40_Re = out_results_40_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_40_Im = out_results_40_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_41_Re = out_results_41_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_41_Im = out_results_41_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_42_Re = out_results_42_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_42_Im = out_results_42_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_43_Re = out_results_43_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_43_Im = out_results_43_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_44_Re = out_results_44_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_44_Im = out_results_44_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_45_Re = out_results_45_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_45_Im = out_results_45_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_46_Re = out_results_46_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_46_Im = out_results_46_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_47_Re = out_results_47_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_47_Im = out_results_47_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_48_Re = out_results_48_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_48_Im = out_results_48_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_49_Re = out_results_49_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_49_Im = out_results_49_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_50_Re = out_results_50_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_50_Im = out_results_50_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_51_Re = out_results_51_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_51_Im = out_results_51_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_52_Re = out_results_52_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_52_Im = out_results_52_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_53_Re = out_results_53_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_53_Im = out_results_53_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_54_Re = out_results_54_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_54_Im = out_results_54_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_55_Re = out_results_55_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_55_Im = out_results_55_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_56_Re = out_results_56_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_56_Im = out_results_56_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_57_Re = out_results_57_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_57_Im = out_results_57_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_58_Re = out_results_58_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_58_Im = out_results_58_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_59_Re = out_results_59_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_59_Im = out_results_59_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_60_Re = out_results_60_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_60_Im = out_results_60_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_61_Re = out_results_61_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_61_Im = out_results_61_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_62_Re = out_results_62_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_62_Im = out_results_62_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_63_Re = out_results_63_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_63_Im = out_results_63_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_64_Re = out_results_64_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_64_Im = out_results_64_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_65_Re = out_results_65_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_65_Im = out_results_65_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_66_Re = out_results_66_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_66_Im = out_results_66_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_67_Re = out_results_67_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_67_Im = out_results_67_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_68_Re = out_results_68_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_68_Im = out_results_68_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_69_Re = out_results_69_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_69_Im = out_results_69_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_70_Re = out_results_70_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_70_Im = out_results_70_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_71_Re = out_results_71_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_71_Im = out_results_71_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_72_Re = out_results_72_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_72_Im = out_results_72_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_73_Re = out_results_73_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_73_Im = out_results_73_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_74_Re = out_results_74_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_74_Im = out_results_74_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_75_Re = out_results_75_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_75_Im = out_results_75_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_76_Re = out_results_76_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_76_Im = out_results_76_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_77_Re = out_results_77_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_77_Im = out_results_77_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_78_Re = out_results_78_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_78_Im = out_results_78_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_79_Re = out_results_79_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_79_Im = out_results_79_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_80_Re = out_results_80_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_80_Im = out_results_80_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_81_Re = out_results_81_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_81_Im = out_results_81_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_82_Re = out_results_82_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_82_Im = out_results_82_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_83_Re = out_results_83_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_83_Im = out_results_83_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_84_Re = out_results_84_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_84_Im = out_results_84_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_85_Re = out_results_85_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_85_Im = out_results_85_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_86_Re = out_results_86_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_86_Im = out_results_86_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_87_Re = out_results_87_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_87_Im = out_results_87_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_88_Re = out_results_88_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_88_Im = out_results_88_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_89_Re = out_results_89_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_89_Im = out_results_89_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_90_Re = out_results_90_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_90_Im = out_results_90_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_91_Re = out_results_91_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_91_Im = out_results_91_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_92_Re = out_results_92_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_92_Im = out_results_92_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_93_Re = out_results_93_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_93_Im = out_results_93_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_94_Re = out_results_94_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_94_Im = out_results_94_Im; // @[FFTDesigns.scala 3474:12]
  assign io_out_95_Re = out_results_95_Re; // @[FFTDesigns.scala 3474:12]
  assign io_out_95_Im = out_results_95_Im; // @[FFTDesigns.scala 3474:12]
  assign FFT_sr_v2_nrv_clock = clock;
  assign FFT_sr_v2_nrv_reset = reset;
  assign FFT_sr_v2_nrv_io_in_0_Re = PermutationsBasic_io_out_0_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_io_in_0_Im = PermutationsBasic_io_out_0_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_io_in_1_Re = PermutationsBasic_io_out_1_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_io_in_1_Im = PermutationsBasic_io_out_1_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_io_in_2_Re = PermutationsBasic_io_out_2_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_io_in_2_Im = PermutationsBasic_io_out_2_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_1_clock = clock;
  assign FFT_sr_v2_nrv_1_reset = reset;
  assign FFT_sr_v2_nrv_1_io_in_0_Re = PermutationsBasic_io_out_3_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_1_io_in_0_Im = PermutationsBasic_io_out_3_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_1_io_in_1_Re = PermutationsBasic_io_out_4_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_1_io_in_1_Im = PermutationsBasic_io_out_4_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_1_io_in_2_Re = PermutationsBasic_io_out_5_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_1_io_in_2_Im = PermutationsBasic_io_out_5_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_2_clock = clock;
  assign FFT_sr_v2_nrv_2_reset = reset;
  assign FFT_sr_v2_nrv_2_io_in_0_Re = PermutationsBasic_io_out_6_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_2_io_in_0_Im = PermutationsBasic_io_out_6_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_2_io_in_1_Re = PermutationsBasic_io_out_7_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_2_io_in_1_Im = PermutationsBasic_io_out_7_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_2_io_in_2_Re = PermutationsBasic_io_out_8_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_2_io_in_2_Im = PermutationsBasic_io_out_8_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_3_clock = clock;
  assign FFT_sr_v2_nrv_3_reset = reset;
  assign FFT_sr_v2_nrv_3_io_in_0_Re = PermutationsBasic_io_out_9_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_3_io_in_0_Im = PermutationsBasic_io_out_9_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_3_io_in_1_Re = PermutationsBasic_io_out_10_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_3_io_in_1_Im = PermutationsBasic_io_out_10_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_3_io_in_2_Re = PermutationsBasic_io_out_11_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_3_io_in_2_Im = PermutationsBasic_io_out_11_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_4_clock = clock;
  assign FFT_sr_v2_nrv_4_reset = reset;
  assign FFT_sr_v2_nrv_4_io_in_0_Re = PermutationsBasic_io_out_12_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_4_io_in_0_Im = PermutationsBasic_io_out_12_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_4_io_in_1_Re = PermutationsBasic_io_out_13_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_4_io_in_1_Im = PermutationsBasic_io_out_13_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_4_io_in_2_Re = PermutationsBasic_io_out_14_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_4_io_in_2_Im = PermutationsBasic_io_out_14_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_5_clock = clock;
  assign FFT_sr_v2_nrv_5_reset = reset;
  assign FFT_sr_v2_nrv_5_io_in_0_Re = PermutationsBasic_io_out_15_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_5_io_in_0_Im = PermutationsBasic_io_out_15_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_5_io_in_1_Re = PermutationsBasic_io_out_16_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_5_io_in_1_Im = PermutationsBasic_io_out_16_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_5_io_in_2_Re = PermutationsBasic_io_out_17_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_5_io_in_2_Im = PermutationsBasic_io_out_17_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_6_clock = clock;
  assign FFT_sr_v2_nrv_6_reset = reset;
  assign FFT_sr_v2_nrv_6_io_in_0_Re = PermutationsBasic_io_out_18_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_6_io_in_0_Im = PermutationsBasic_io_out_18_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_6_io_in_1_Re = PermutationsBasic_io_out_19_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_6_io_in_1_Im = PermutationsBasic_io_out_19_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_6_io_in_2_Re = PermutationsBasic_io_out_20_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_6_io_in_2_Im = PermutationsBasic_io_out_20_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_7_clock = clock;
  assign FFT_sr_v2_nrv_7_reset = reset;
  assign FFT_sr_v2_nrv_7_io_in_0_Re = PermutationsBasic_io_out_21_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_7_io_in_0_Im = PermutationsBasic_io_out_21_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_7_io_in_1_Re = PermutationsBasic_io_out_22_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_7_io_in_1_Im = PermutationsBasic_io_out_22_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_7_io_in_2_Re = PermutationsBasic_io_out_23_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_7_io_in_2_Im = PermutationsBasic_io_out_23_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_8_clock = clock;
  assign FFT_sr_v2_nrv_8_reset = reset;
  assign FFT_sr_v2_nrv_8_io_in_0_Re = PermutationsBasic_io_out_24_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_8_io_in_0_Im = PermutationsBasic_io_out_24_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_8_io_in_1_Re = PermutationsBasic_io_out_25_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_8_io_in_1_Im = PermutationsBasic_io_out_25_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_8_io_in_2_Re = PermutationsBasic_io_out_26_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_8_io_in_2_Im = PermutationsBasic_io_out_26_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_9_clock = clock;
  assign FFT_sr_v2_nrv_9_reset = reset;
  assign FFT_sr_v2_nrv_9_io_in_0_Re = PermutationsBasic_io_out_27_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_9_io_in_0_Im = PermutationsBasic_io_out_27_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_9_io_in_1_Re = PermutationsBasic_io_out_28_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_9_io_in_1_Im = PermutationsBasic_io_out_28_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_9_io_in_2_Re = PermutationsBasic_io_out_29_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_9_io_in_2_Im = PermutationsBasic_io_out_29_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_10_clock = clock;
  assign FFT_sr_v2_nrv_10_reset = reset;
  assign FFT_sr_v2_nrv_10_io_in_0_Re = PermutationsBasic_io_out_30_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_10_io_in_0_Im = PermutationsBasic_io_out_30_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_10_io_in_1_Re = PermutationsBasic_io_out_31_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_10_io_in_1_Im = PermutationsBasic_io_out_31_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_10_io_in_2_Re = PermutationsBasic_io_out_32_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_10_io_in_2_Im = PermutationsBasic_io_out_32_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_11_clock = clock;
  assign FFT_sr_v2_nrv_11_reset = reset;
  assign FFT_sr_v2_nrv_11_io_in_0_Re = PermutationsBasic_io_out_33_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_11_io_in_0_Im = PermutationsBasic_io_out_33_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_11_io_in_1_Re = PermutationsBasic_io_out_34_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_11_io_in_1_Im = PermutationsBasic_io_out_34_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_11_io_in_2_Re = PermutationsBasic_io_out_35_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_11_io_in_2_Im = PermutationsBasic_io_out_35_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_12_clock = clock;
  assign FFT_sr_v2_nrv_12_reset = reset;
  assign FFT_sr_v2_nrv_12_io_in_0_Re = PermutationsBasic_io_out_36_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_12_io_in_0_Im = PermutationsBasic_io_out_36_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_12_io_in_1_Re = PermutationsBasic_io_out_37_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_12_io_in_1_Im = PermutationsBasic_io_out_37_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_12_io_in_2_Re = PermutationsBasic_io_out_38_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_12_io_in_2_Im = PermutationsBasic_io_out_38_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_13_clock = clock;
  assign FFT_sr_v2_nrv_13_reset = reset;
  assign FFT_sr_v2_nrv_13_io_in_0_Re = PermutationsBasic_io_out_39_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_13_io_in_0_Im = PermutationsBasic_io_out_39_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_13_io_in_1_Re = PermutationsBasic_io_out_40_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_13_io_in_1_Im = PermutationsBasic_io_out_40_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_13_io_in_2_Re = PermutationsBasic_io_out_41_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_13_io_in_2_Im = PermutationsBasic_io_out_41_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_14_clock = clock;
  assign FFT_sr_v2_nrv_14_reset = reset;
  assign FFT_sr_v2_nrv_14_io_in_0_Re = PermutationsBasic_io_out_42_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_14_io_in_0_Im = PermutationsBasic_io_out_42_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_14_io_in_1_Re = PermutationsBasic_io_out_43_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_14_io_in_1_Im = PermutationsBasic_io_out_43_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_14_io_in_2_Re = PermutationsBasic_io_out_44_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_14_io_in_2_Im = PermutationsBasic_io_out_44_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_15_clock = clock;
  assign FFT_sr_v2_nrv_15_reset = reset;
  assign FFT_sr_v2_nrv_15_io_in_0_Re = PermutationsBasic_io_out_45_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_15_io_in_0_Im = PermutationsBasic_io_out_45_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_15_io_in_1_Re = PermutationsBasic_io_out_46_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_15_io_in_1_Im = PermutationsBasic_io_out_46_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_15_io_in_2_Re = PermutationsBasic_io_out_47_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_15_io_in_2_Im = PermutationsBasic_io_out_47_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_16_clock = clock;
  assign FFT_sr_v2_nrv_16_reset = reset;
  assign FFT_sr_v2_nrv_16_io_in_0_Re = PermutationsBasic_io_out_48_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_16_io_in_0_Im = PermutationsBasic_io_out_48_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_16_io_in_1_Re = PermutationsBasic_io_out_49_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_16_io_in_1_Im = PermutationsBasic_io_out_49_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_16_io_in_2_Re = PermutationsBasic_io_out_50_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_16_io_in_2_Im = PermutationsBasic_io_out_50_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_17_clock = clock;
  assign FFT_sr_v2_nrv_17_reset = reset;
  assign FFT_sr_v2_nrv_17_io_in_0_Re = PermutationsBasic_io_out_51_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_17_io_in_0_Im = PermutationsBasic_io_out_51_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_17_io_in_1_Re = PermutationsBasic_io_out_52_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_17_io_in_1_Im = PermutationsBasic_io_out_52_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_17_io_in_2_Re = PermutationsBasic_io_out_53_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_17_io_in_2_Im = PermutationsBasic_io_out_53_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_18_clock = clock;
  assign FFT_sr_v2_nrv_18_reset = reset;
  assign FFT_sr_v2_nrv_18_io_in_0_Re = PermutationsBasic_io_out_54_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_18_io_in_0_Im = PermutationsBasic_io_out_54_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_18_io_in_1_Re = PermutationsBasic_io_out_55_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_18_io_in_1_Im = PermutationsBasic_io_out_55_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_18_io_in_2_Re = PermutationsBasic_io_out_56_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_18_io_in_2_Im = PermutationsBasic_io_out_56_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_19_clock = clock;
  assign FFT_sr_v2_nrv_19_reset = reset;
  assign FFT_sr_v2_nrv_19_io_in_0_Re = PermutationsBasic_io_out_57_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_19_io_in_0_Im = PermutationsBasic_io_out_57_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_19_io_in_1_Re = PermutationsBasic_io_out_58_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_19_io_in_1_Im = PermutationsBasic_io_out_58_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_19_io_in_2_Re = PermutationsBasic_io_out_59_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_19_io_in_2_Im = PermutationsBasic_io_out_59_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_20_clock = clock;
  assign FFT_sr_v2_nrv_20_reset = reset;
  assign FFT_sr_v2_nrv_20_io_in_0_Re = PermutationsBasic_io_out_60_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_20_io_in_0_Im = PermutationsBasic_io_out_60_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_20_io_in_1_Re = PermutationsBasic_io_out_61_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_20_io_in_1_Im = PermutationsBasic_io_out_61_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_20_io_in_2_Re = PermutationsBasic_io_out_62_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_20_io_in_2_Im = PermutationsBasic_io_out_62_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_21_clock = clock;
  assign FFT_sr_v2_nrv_21_reset = reset;
  assign FFT_sr_v2_nrv_21_io_in_0_Re = PermutationsBasic_io_out_63_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_21_io_in_0_Im = PermutationsBasic_io_out_63_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_21_io_in_1_Re = PermutationsBasic_io_out_64_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_21_io_in_1_Im = PermutationsBasic_io_out_64_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_21_io_in_2_Re = PermutationsBasic_io_out_65_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_21_io_in_2_Im = PermutationsBasic_io_out_65_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_22_clock = clock;
  assign FFT_sr_v2_nrv_22_reset = reset;
  assign FFT_sr_v2_nrv_22_io_in_0_Re = PermutationsBasic_io_out_66_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_22_io_in_0_Im = PermutationsBasic_io_out_66_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_22_io_in_1_Re = PermutationsBasic_io_out_67_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_22_io_in_1_Im = PermutationsBasic_io_out_67_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_22_io_in_2_Re = PermutationsBasic_io_out_68_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_22_io_in_2_Im = PermutationsBasic_io_out_68_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_23_clock = clock;
  assign FFT_sr_v2_nrv_23_reset = reset;
  assign FFT_sr_v2_nrv_23_io_in_0_Re = PermutationsBasic_io_out_69_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_23_io_in_0_Im = PermutationsBasic_io_out_69_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_23_io_in_1_Re = PermutationsBasic_io_out_70_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_23_io_in_1_Im = PermutationsBasic_io_out_70_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_23_io_in_2_Re = PermutationsBasic_io_out_71_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_23_io_in_2_Im = PermutationsBasic_io_out_71_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_24_clock = clock;
  assign FFT_sr_v2_nrv_24_reset = reset;
  assign FFT_sr_v2_nrv_24_io_in_0_Re = PermutationsBasic_io_out_72_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_24_io_in_0_Im = PermutationsBasic_io_out_72_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_24_io_in_1_Re = PermutationsBasic_io_out_73_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_24_io_in_1_Im = PermutationsBasic_io_out_73_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_24_io_in_2_Re = PermutationsBasic_io_out_74_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_24_io_in_2_Im = PermutationsBasic_io_out_74_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_25_clock = clock;
  assign FFT_sr_v2_nrv_25_reset = reset;
  assign FFT_sr_v2_nrv_25_io_in_0_Re = PermutationsBasic_io_out_75_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_25_io_in_0_Im = PermutationsBasic_io_out_75_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_25_io_in_1_Re = PermutationsBasic_io_out_76_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_25_io_in_1_Im = PermutationsBasic_io_out_76_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_25_io_in_2_Re = PermutationsBasic_io_out_77_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_25_io_in_2_Im = PermutationsBasic_io_out_77_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_26_clock = clock;
  assign FFT_sr_v2_nrv_26_reset = reset;
  assign FFT_sr_v2_nrv_26_io_in_0_Re = PermutationsBasic_io_out_78_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_26_io_in_0_Im = PermutationsBasic_io_out_78_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_26_io_in_1_Re = PermutationsBasic_io_out_79_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_26_io_in_1_Im = PermutationsBasic_io_out_79_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_26_io_in_2_Re = PermutationsBasic_io_out_80_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_26_io_in_2_Im = PermutationsBasic_io_out_80_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_27_clock = clock;
  assign FFT_sr_v2_nrv_27_reset = reset;
  assign FFT_sr_v2_nrv_27_io_in_0_Re = PermutationsBasic_io_out_81_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_27_io_in_0_Im = PermutationsBasic_io_out_81_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_27_io_in_1_Re = PermutationsBasic_io_out_82_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_27_io_in_1_Im = PermutationsBasic_io_out_82_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_27_io_in_2_Re = PermutationsBasic_io_out_83_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_27_io_in_2_Im = PermutationsBasic_io_out_83_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_28_clock = clock;
  assign FFT_sr_v2_nrv_28_reset = reset;
  assign FFT_sr_v2_nrv_28_io_in_0_Re = PermutationsBasic_io_out_84_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_28_io_in_0_Im = PermutationsBasic_io_out_84_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_28_io_in_1_Re = PermutationsBasic_io_out_85_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_28_io_in_1_Im = PermutationsBasic_io_out_85_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_28_io_in_2_Re = PermutationsBasic_io_out_86_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_28_io_in_2_Im = PermutationsBasic_io_out_86_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_29_clock = clock;
  assign FFT_sr_v2_nrv_29_reset = reset;
  assign FFT_sr_v2_nrv_29_io_in_0_Re = PermutationsBasic_io_out_87_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_29_io_in_0_Im = PermutationsBasic_io_out_87_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_29_io_in_1_Re = PermutationsBasic_io_out_88_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_29_io_in_1_Im = PermutationsBasic_io_out_88_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_29_io_in_2_Re = PermutationsBasic_io_out_89_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_29_io_in_2_Im = PermutationsBasic_io_out_89_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_30_clock = clock;
  assign FFT_sr_v2_nrv_30_reset = reset;
  assign FFT_sr_v2_nrv_30_io_in_0_Re = PermutationsBasic_io_out_90_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_30_io_in_0_Im = PermutationsBasic_io_out_90_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_30_io_in_1_Re = PermutationsBasic_io_out_91_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_30_io_in_1_Im = PermutationsBasic_io_out_91_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_30_io_in_2_Re = PermutationsBasic_io_out_92_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_30_io_in_2_Im = PermutationsBasic_io_out_92_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_31_clock = clock;
  assign FFT_sr_v2_nrv_31_reset = reset;
  assign FFT_sr_v2_nrv_31_io_in_0_Re = PermutationsBasic_io_out_93_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_31_io_in_0_Im = PermutationsBasic_io_out_93_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_31_io_in_1_Re = PermutationsBasic_io_out_94_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_31_io_in_1_Im = PermutationsBasic_io_out_94_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_31_io_in_2_Re = PermutationsBasic_io_out_95_Re; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_31_io_in_2_Im = PermutationsBasic_io_out_95_Im; // @[FFTDesigns.scala 3477:32]
  assign FFT_sr_v2_nrv_32_clock = clock;
  assign FFT_sr_v2_nrv_32_reset = reset;
  assign FFT_sr_v2_nrv_32_io_in_0_Re = TwiddleFactors_mr_io_out_0_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_0_Im = TwiddleFactors_mr_io_out_0_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_1_Re = TwiddleFactors_mr_io_out_1_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_1_Im = TwiddleFactors_mr_io_out_1_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_2_Re = TwiddleFactors_mr_io_out_2_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_2_Im = TwiddleFactors_mr_io_out_2_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_3_Re = TwiddleFactors_mr_io_out_3_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_3_Im = TwiddleFactors_mr_io_out_3_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_4_Re = TwiddleFactors_mr_io_out_4_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_4_Im = TwiddleFactors_mr_io_out_4_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_5_Re = TwiddleFactors_mr_io_out_5_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_5_Im = TwiddleFactors_mr_io_out_5_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_6_Re = TwiddleFactors_mr_io_out_6_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_6_Im = TwiddleFactors_mr_io_out_6_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_7_Re = TwiddleFactors_mr_io_out_7_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_7_Im = TwiddleFactors_mr_io_out_7_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_8_Re = TwiddleFactors_mr_io_out_8_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_8_Im = TwiddleFactors_mr_io_out_8_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_9_Re = TwiddleFactors_mr_io_out_9_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_9_Im = TwiddleFactors_mr_io_out_9_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_10_Re = TwiddleFactors_mr_io_out_10_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_10_Im = TwiddleFactors_mr_io_out_10_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_11_Re = TwiddleFactors_mr_io_out_11_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_11_Im = TwiddleFactors_mr_io_out_11_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_12_Re = TwiddleFactors_mr_io_out_12_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_12_Im = TwiddleFactors_mr_io_out_12_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_13_Re = TwiddleFactors_mr_io_out_13_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_13_Im = TwiddleFactors_mr_io_out_13_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_14_Re = TwiddleFactors_mr_io_out_14_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_14_Im = TwiddleFactors_mr_io_out_14_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_15_Re = TwiddleFactors_mr_io_out_15_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_15_Im = TwiddleFactors_mr_io_out_15_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_16_Re = TwiddleFactors_mr_io_out_16_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_16_Im = TwiddleFactors_mr_io_out_16_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_17_Re = TwiddleFactors_mr_io_out_17_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_17_Im = TwiddleFactors_mr_io_out_17_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_18_Re = TwiddleFactors_mr_io_out_18_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_18_Im = TwiddleFactors_mr_io_out_18_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_19_Re = TwiddleFactors_mr_io_out_19_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_19_Im = TwiddleFactors_mr_io_out_19_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_20_Re = TwiddleFactors_mr_io_out_20_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_20_Im = TwiddleFactors_mr_io_out_20_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_21_Re = TwiddleFactors_mr_io_out_21_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_21_Im = TwiddleFactors_mr_io_out_21_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_22_Re = TwiddleFactors_mr_io_out_22_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_22_Im = TwiddleFactors_mr_io_out_22_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_23_Re = TwiddleFactors_mr_io_out_23_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_23_Im = TwiddleFactors_mr_io_out_23_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_24_Re = TwiddleFactors_mr_io_out_24_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_24_Im = TwiddleFactors_mr_io_out_24_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_25_Re = TwiddleFactors_mr_io_out_25_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_25_Im = TwiddleFactors_mr_io_out_25_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_26_Re = TwiddleFactors_mr_io_out_26_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_26_Im = TwiddleFactors_mr_io_out_26_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_27_Re = TwiddleFactors_mr_io_out_27_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_27_Im = TwiddleFactors_mr_io_out_27_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_28_Re = TwiddleFactors_mr_io_out_28_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_28_Im = TwiddleFactors_mr_io_out_28_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_29_Re = TwiddleFactors_mr_io_out_29_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_29_Im = TwiddleFactors_mr_io_out_29_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_30_Re = TwiddleFactors_mr_io_out_30_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_30_Im = TwiddleFactors_mr_io_out_30_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_31_Re = TwiddleFactors_mr_io_out_31_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_32_io_in_31_Im = TwiddleFactors_mr_io_out_31_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_clock = clock;
  assign FFT_sr_v2_nrv_33_reset = reset;
  assign FFT_sr_v2_nrv_33_io_in_0_Re = TwiddleFactors_mr_io_out_32_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_0_Im = TwiddleFactors_mr_io_out_32_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_1_Re = TwiddleFactors_mr_io_out_33_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_1_Im = TwiddleFactors_mr_io_out_33_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_2_Re = TwiddleFactors_mr_io_out_34_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_2_Im = TwiddleFactors_mr_io_out_34_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_3_Re = TwiddleFactors_mr_io_out_35_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_3_Im = TwiddleFactors_mr_io_out_35_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_4_Re = TwiddleFactors_mr_io_out_36_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_4_Im = TwiddleFactors_mr_io_out_36_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_5_Re = TwiddleFactors_mr_io_out_37_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_5_Im = TwiddleFactors_mr_io_out_37_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_6_Re = TwiddleFactors_mr_io_out_38_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_6_Im = TwiddleFactors_mr_io_out_38_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_7_Re = TwiddleFactors_mr_io_out_39_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_7_Im = TwiddleFactors_mr_io_out_39_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_8_Re = TwiddleFactors_mr_io_out_40_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_8_Im = TwiddleFactors_mr_io_out_40_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_9_Re = TwiddleFactors_mr_io_out_41_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_9_Im = TwiddleFactors_mr_io_out_41_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_10_Re = TwiddleFactors_mr_io_out_42_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_10_Im = TwiddleFactors_mr_io_out_42_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_11_Re = TwiddleFactors_mr_io_out_43_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_11_Im = TwiddleFactors_mr_io_out_43_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_12_Re = TwiddleFactors_mr_io_out_44_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_12_Im = TwiddleFactors_mr_io_out_44_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_13_Re = TwiddleFactors_mr_io_out_45_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_13_Im = TwiddleFactors_mr_io_out_45_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_14_Re = TwiddleFactors_mr_io_out_46_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_14_Im = TwiddleFactors_mr_io_out_46_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_15_Re = TwiddleFactors_mr_io_out_47_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_15_Im = TwiddleFactors_mr_io_out_47_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_16_Re = TwiddleFactors_mr_io_out_48_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_16_Im = TwiddleFactors_mr_io_out_48_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_17_Re = TwiddleFactors_mr_io_out_49_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_17_Im = TwiddleFactors_mr_io_out_49_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_18_Re = TwiddleFactors_mr_io_out_50_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_18_Im = TwiddleFactors_mr_io_out_50_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_19_Re = TwiddleFactors_mr_io_out_51_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_19_Im = TwiddleFactors_mr_io_out_51_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_20_Re = TwiddleFactors_mr_io_out_52_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_20_Im = TwiddleFactors_mr_io_out_52_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_21_Re = TwiddleFactors_mr_io_out_53_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_21_Im = TwiddleFactors_mr_io_out_53_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_22_Re = TwiddleFactors_mr_io_out_54_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_22_Im = TwiddleFactors_mr_io_out_54_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_23_Re = TwiddleFactors_mr_io_out_55_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_23_Im = TwiddleFactors_mr_io_out_55_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_24_Re = TwiddleFactors_mr_io_out_56_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_24_Im = TwiddleFactors_mr_io_out_56_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_25_Re = TwiddleFactors_mr_io_out_57_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_25_Im = TwiddleFactors_mr_io_out_57_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_26_Re = TwiddleFactors_mr_io_out_58_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_26_Im = TwiddleFactors_mr_io_out_58_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_27_Re = TwiddleFactors_mr_io_out_59_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_27_Im = TwiddleFactors_mr_io_out_59_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_28_Re = TwiddleFactors_mr_io_out_60_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_28_Im = TwiddleFactors_mr_io_out_60_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_29_Re = TwiddleFactors_mr_io_out_61_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_29_Im = TwiddleFactors_mr_io_out_61_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_30_Re = TwiddleFactors_mr_io_out_62_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_30_Im = TwiddleFactors_mr_io_out_62_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_31_Re = TwiddleFactors_mr_io_out_63_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_33_io_in_31_Im = TwiddleFactors_mr_io_out_63_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_clock = clock;
  assign FFT_sr_v2_nrv_34_reset = reset;
  assign FFT_sr_v2_nrv_34_io_in_0_Re = TwiddleFactors_mr_io_out_64_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_0_Im = TwiddleFactors_mr_io_out_64_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_1_Re = TwiddleFactors_mr_io_out_65_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_1_Im = TwiddleFactors_mr_io_out_65_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_2_Re = TwiddleFactors_mr_io_out_66_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_2_Im = TwiddleFactors_mr_io_out_66_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_3_Re = TwiddleFactors_mr_io_out_67_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_3_Im = TwiddleFactors_mr_io_out_67_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_4_Re = TwiddleFactors_mr_io_out_68_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_4_Im = TwiddleFactors_mr_io_out_68_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_5_Re = TwiddleFactors_mr_io_out_69_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_5_Im = TwiddleFactors_mr_io_out_69_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_6_Re = TwiddleFactors_mr_io_out_70_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_6_Im = TwiddleFactors_mr_io_out_70_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_7_Re = TwiddleFactors_mr_io_out_71_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_7_Im = TwiddleFactors_mr_io_out_71_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_8_Re = TwiddleFactors_mr_io_out_72_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_8_Im = TwiddleFactors_mr_io_out_72_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_9_Re = TwiddleFactors_mr_io_out_73_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_9_Im = TwiddleFactors_mr_io_out_73_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_10_Re = TwiddleFactors_mr_io_out_74_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_10_Im = TwiddleFactors_mr_io_out_74_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_11_Re = TwiddleFactors_mr_io_out_75_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_11_Im = TwiddleFactors_mr_io_out_75_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_12_Re = TwiddleFactors_mr_io_out_76_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_12_Im = TwiddleFactors_mr_io_out_76_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_13_Re = TwiddleFactors_mr_io_out_77_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_13_Im = TwiddleFactors_mr_io_out_77_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_14_Re = TwiddleFactors_mr_io_out_78_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_14_Im = TwiddleFactors_mr_io_out_78_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_15_Re = TwiddleFactors_mr_io_out_79_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_15_Im = TwiddleFactors_mr_io_out_79_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_16_Re = TwiddleFactors_mr_io_out_80_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_16_Im = TwiddleFactors_mr_io_out_80_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_17_Re = TwiddleFactors_mr_io_out_81_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_17_Im = TwiddleFactors_mr_io_out_81_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_18_Re = TwiddleFactors_mr_io_out_82_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_18_Im = TwiddleFactors_mr_io_out_82_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_19_Re = TwiddleFactors_mr_io_out_83_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_19_Im = TwiddleFactors_mr_io_out_83_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_20_Re = TwiddleFactors_mr_io_out_84_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_20_Im = TwiddleFactors_mr_io_out_84_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_21_Re = TwiddleFactors_mr_io_out_85_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_21_Im = TwiddleFactors_mr_io_out_85_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_22_Re = TwiddleFactors_mr_io_out_86_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_22_Im = TwiddleFactors_mr_io_out_86_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_23_Re = TwiddleFactors_mr_io_out_87_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_23_Im = TwiddleFactors_mr_io_out_87_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_24_Re = TwiddleFactors_mr_io_out_88_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_24_Im = TwiddleFactors_mr_io_out_88_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_25_Re = TwiddleFactors_mr_io_out_89_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_25_Im = TwiddleFactors_mr_io_out_89_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_26_Re = TwiddleFactors_mr_io_out_90_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_26_Im = TwiddleFactors_mr_io_out_90_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_27_Re = TwiddleFactors_mr_io_out_91_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_27_Im = TwiddleFactors_mr_io_out_91_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_28_Re = TwiddleFactors_mr_io_out_92_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_28_Im = TwiddleFactors_mr_io_out_92_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_29_Re = TwiddleFactors_mr_io_out_93_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_29_Im = TwiddleFactors_mr_io_out_93_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_30_Re = TwiddleFactors_mr_io_out_94_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_30_Im = TwiddleFactors_mr_io_out_94_Im; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_31_Re = TwiddleFactors_mr_io_out_95_Re; // @[FFTDesigns.scala 3479:32]
  assign FFT_sr_v2_nrv_34_io_in_31_Im = TwiddleFactors_mr_io_out_95_Im; // @[FFTDesigns.scala 3479:32]
  assign PermutationsBasic_io_in_0_Re = io_in_ready ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_0_Im = io_in_ready ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_1_Re = io_in_ready ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_1_Im = io_in_ready ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_2_Re = io_in_ready ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_2_Im = io_in_ready ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_3_Re = io_in_ready ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_3_Im = io_in_ready ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_4_Re = io_in_ready ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_4_Im = io_in_ready ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_5_Re = io_in_ready ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_5_Im = io_in_ready ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_6_Re = io_in_ready ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_6_Im = io_in_ready ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_7_Re = io_in_ready ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_7_Im = io_in_ready ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_8_Re = io_in_ready ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_8_Im = io_in_ready ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_9_Re = io_in_ready ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_9_Im = io_in_ready ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_10_Re = io_in_ready ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_10_Im = io_in_ready ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_11_Re = io_in_ready ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_11_Im = io_in_ready ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_12_Re = io_in_ready ? io_in_12_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_12_Im = io_in_ready ? io_in_12_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_13_Re = io_in_ready ? io_in_13_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_13_Im = io_in_ready ? io_in_13_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_14_Re = io_in_ready ? io_in_14_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_14_Im = io_in_ready ? io_in_14_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_15_Re = io_in_ready ? io_in_15_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_15_Im = io_in_ready ? io_in_15_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_16_Re = io_in_ready ? io_in_16_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_16_Im = io_in_ready ? io_in_16_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_17_Re = io_in_ready ? io_in_17_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_17_Im = io_in_ready ? io_in_17_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_18_Re = io_in_ready ? io_in_18_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_18_Im = io_in_ready ? io_in_18_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_19_Re = io_in_ready ? io_in_19_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_19_Im = io_in_ready ? io_in_19_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_20_Re = io_in_ready ? io_in_20_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_20_Im = io_in_ready ? io_in_20_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_21_Re = io_in_ready ? io_in_21_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_21_Im = io_in_ready ? io_in_21_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_22_Re = io_in_ready ? io_in_22_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_22_Im = io_in_ready ? io_in_22_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_23_Re = io_in_ready ? io_in_23_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_23_Im = io_in_ready ? io_in_23_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_24_Re = io_in_ready ? io_in_24_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_24_Im = io_in_ready ? io_in_24_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_25_Re = io_in_ready ? io_in_25_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_25_Im = io_in_ready ? io_in_25_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_26_Re = io_in_ready ? io_in_26_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_26_Im = io_in_ready ? io_in_26_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_27_Re = io_in_ready ? io_in_27_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_27_Im = io_in_ready ? io_in_27_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_28_Re = io_in_ready ? io_in_28_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_28_Im = io_in_ready ? io_in_28_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_29_Re = io_in_ready ? io_in_29_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_29_Im = io_in_ready ? io_in_29_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_30_Re = io_in_ready ? io_in_30_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_30_Im = io_in_ready ? io_in_30_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_31_Re = io_in_ready ? io_in_31_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_31_Im = io_in_ready ? io_in_31_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_32_Re = io_in_ready ? io_in_32_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_32_Im = io_in_ready ? io_in_32_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_33_Re = io_in_ready ? io_in_33_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_33_Im = io_in_ready ? io_in_33_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_34_Re = io_in_ready ? io_in_34_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_34_Im = io_in_ready ? io_in_34_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_35_Re = io_in_ready ? io_in_35_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_35_Im = io_in_ready ? io_in_35_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_36_Re = io_in_ready ? io_in_36_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_36_Im = io_in_ready ? io_in_36_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_37_Re = io_in_ready ? io_in_37_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_37_Im = io_in_ready ? io_in_37_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_38_Re = io_in_ready ? io_in_38_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_38_Im = io_in_ready ? io_in_38_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_39_Re = io_in_ready ? io_in_39_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_39_Im = io_in_ready ? io_in_39_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_40_Re = io_in_ready ? io_in_40_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_40_Im = io_in_ready ? io_in_40_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_41_Re = io_in_ready ? io_in_41_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_41_Im = io_in_ready ? io_in_41_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_42_Re = io_in_ready ? io_in_42_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_42_Im = io_in_ready ? io_in_42_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_43_Re = io_in_ready ? io_in_43_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_43_Im = io_in_ready ? io_in_43_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_44_Re = io_in_ready ? io_in_44_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_44_Im = io_in_ready ? io_in_44_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_45_Re = io_in_ready ? io_in_45_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_45_Im = io_in_ready ? io_in_45_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_46_Re = io_in_ready ? io_in_46_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_46_Im = io_in_ready ? io_in_46_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_47_Re = io_in_ready ? io_in_47_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_47_Im = io_in_ready ? io_in_47_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_48_Re = io_in_ready ? io_in_48_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_48_Im = io_in_ready ? io_in_48_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_49_Re = io_in_ready ? io_in_49_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_49_Im = io_in_ready ? io_in_49_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_50_Re = io_in_ready ? io_in_50_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_50_Im = io_in_ready ? io_in_50_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_51_Re = io_in_ready ? io_in_51_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_51_Im = io_in_ready ? io_in_51_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_52_Re = io_in_ready ? io_in_52_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_52_Im = io_in_ready ? io_in_52_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_53_Re = io_in_ready ? io_in_53_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_53_Im = io_in_ready ? io_in_53_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_54_Re = io_in_ready ? io_in_54_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_54_Im = io_in_ready ? io_in_54_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_55_Re = io_in_ready ? io_in_55_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_55_Im = io_in_ready ? io_in_55_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_56_Re = io_in_ready ? io_in_56_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_56_Im = io_in_ready ? io_in_56_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_57_Re = io_in_ready ? io_in_57_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_57_Im = io_in_ready ? io_in_57_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_58_Re = io_in_ready ? io_in_58_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_58_Im = io_in_ready ? io_in_58_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_59_Re = io_in_ready ? io_in_59_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_59_Im = io_in_ready ? io_in_59_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_60_Re = io_in_ready ? io_in_60_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_60_Im = io_in_ready ? io_in_60_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_61_Re = io_in_ready ? io_in_61_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_61_Im = io_in_ready ? io_in_61_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_62_Re = io_in_ready ? io_in_62_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_62_Im = io_in_ready ? io_in_62_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_63_Re = io_in_ready ? io_in_63_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_63_Im = io_in_ready ? io_in_63_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_64_Re = io_in_ready ? io_in_64_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_64_Im = io_in_ready ? io_in_64_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_65_Re = io_in_ready ? io_in_65_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_65_Im = io_in_ready ? io_in_65_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_66_Re = io_in_ready ? io_in_66_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_66_Im = io_in_ready ? io_in_66_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_67_Re = io_in_ready ? io_in_67_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_67_Im = io_in_ready ? io_in_67_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_68_Re = io_in_ready ? io_in_68_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_68_Im = io_in_ready ? io_in_68_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_69_Re = io_in_ready ? io_in_69_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_69_Im = io_in_ready ? io_in_69_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_70_Re = io_in_ready ? io_in_70_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_70_Im = io_in_ready ? io_in_70_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_71_Re = io_in_ready ? io_in_71_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_71_Im = io_in_ready ? io_in_71_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_72_Re = io_in_ready ? io_in_72_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_72_Im = io_in_ready ? io_in_72_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_73_Re = io_in_ready ? io_in_73_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_73_Im = io_in_ready ? io_in_73_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_74_Re = io_in_ready ? io_in_74_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_74_Im = io_in_ready ? io_in_74_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_75_Re = io_in_ready ? io_in_75_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_75_Im = io_in_ready ? io_in_75_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_76_Re = io_in_ready ? io_in_76_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_76_Im = io_in_ready ? io_in_76_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_77_Re = io_in_ready ? io_in_77_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_77_Im = io_in_ready ? io_in_77_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_78_Re = io_in_ready ? io_in_78_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_78_Im = io_in_ready ? io_in_78_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_79_Re = io_in_ready ? io_in_79_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_79_Im = io_in_ready ? io_in_79_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_80_Re = io_in_ready ? io_in_80_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_80_Im = io_in_ready ? io_in_80_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_81_Re = io_in_ready ? io_in_81_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_81_Im = io_in_ready ? io_in_81_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_82_Re = io_in_ready ? io_in_82_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_82_Im = io_in_ready ? io_in_82_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_83_Re = io_in_ready ? io_in_83_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_83_Im = io_in_ready ? io_in_83_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_84_Re = io_in_ready ? io_in_84_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_84_Im = io_in_ready ? io_in_84_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_85_Re = io_in_ready ? io_in_85_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_85_Im = io_in_ready ? io_in_85_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_86_Re = io_in_ready ? io_in_86_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_86_Im = io_in_ready ? io_in_86_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_87_Re = io_in_ready ? io_in_87_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_87_Im = io_in_ready ? io_in_87_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_88_Re = io_in_ready ? io_in_88_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_88_Im = io_in_ready ? io_in_88_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_89_Re = io_in_ready ? io_in_89_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_89_Im = io_in_ready ? io_in_89_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_90_Re = io_in_ready ? io_in_90_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_90_Im = io_in_ready ? io_in_90_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_91_Re = io_in_ready ? io_in_91_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_91_Im = io_in_ready ? io_in_91_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_92_Re = io_in_ready ? io_in_92_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_92_Im = io_in_ready ? io_in_92_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_93_Re = io_in_ready ? io_in_93_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_93_Im = io_in_ready ? io_in_93_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_94_Re = io_in_ready ? io_in_94_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_94_Im = io_in_ready ? io_in_94_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_95_Re = io_in_ready ? io_in_95_Re : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_io_in_95_Im = io_in_ready ? io_in_95_Im : 32'h0; // @[FFTDesigns.scala 3455:22 3456:33 3459:38]
  assign PermutationsBasic_1_io_in_0_Re = FFT_sr_v2_nrv_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_0_Im = FFT_sr_v2_nrv_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_1_Re = FFT_sr_v2_nrv_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_1_Im = FFT_sr_v2_nrv_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_2_Re = FFT_sr_v2_nrv_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_2_Im = FFT_sr_v2_nrv_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_3_Re = FFT_sr_v2_nrv_1_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_3_Im = FFT_sr_v2_nrv_1_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_4_Re = FFT_sr_v2_nrv_1_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_4_Im = FFT_sr_v2_nrv_1_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_5_Re = FFT_sr_v2_nrv_1_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_5_Im = FFT_sr_v2_nrv_1_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_6_Re = FFT_sr_v2_nrv_2_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_6_Im = FFT_sr_v2_nrv_2_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_7_Re = FFT_sr_v2_nrv_2_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_7_Im = FFT_sr_v2_nrv_2_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_8_Re = FFT_sr_v2_nrv_2_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_8_Im = FFT_sr_v2_nrv_2_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_9_Re = FFT_sr_v2_nrv_3_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_9_Im = FFT_sr_v2_nrv_3_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_10_Re = FFT_sr_v2_nrv_3_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_10_Im = FFT_sr_v2_nrv_3_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_11_Re = FFT_sr_v2_nrv_3_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_11_Im = FFT_sr_v2_nrv_3_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_12_Re = FFT_sr_v2_nrv_4_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_12_Im = FFT_sr_v2_nrv_4_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_13_Re = FFT_sr_v2_nrv_4_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_13_Im = FFT_sr_v2_nrv_4_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_14_Re = FFT_sr_v2_nrv_4_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_14_Im = FFT_sr_v2_nrv_4_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_15_Re = FFT_sr_v2_nrv_5_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_15_Im = FFT_sr_v2_nrv_5_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_16_Re = FFT_sr_v2_nrv_5_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_16_Im = FFT_sr_v2_nrv_5_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_17_Re = FFT_sr_v2_nrv_5_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_17_Im = FFT_sr_v2_nrv_5_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_18_Re = FFT_sr_v2_nrv_6_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_18_Im = FFT_sr_v2_nrv_6_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_19_Re = FFT_sr_v2_nrv_6_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_19_Im = FFT_sr_v2_nrv_6_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_20_Re = FFT_sr_v2_nrv_6_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_20_Im = FFT_sr_v2_nrv_6_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_21_Re = FFT_sr_v2_nrv_7_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_21_Im = FFT_sr_v2_nrv_7_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_22_Re = FFT_sr_v2_nrv_7_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_22_Im = FFT_sr_v2_nrv_7_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_23_Re = FFT_sr_v2_nrv_7_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_23_Im = FFT_sr_v2_nrv_7_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_24_Re = FFT_sr_v2_nrv_8_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_24_Im = FFT_sr_v2_nrv_8_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_25_Re = FFT_sr_v2_nrv_8_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_25_Im = FFT_sr_v2_nrv_8_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_26_Re = FFT_sr_v2_nrv_8_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_26_Im = FFT_sr_v2_nrv_8_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_27_Re = FFT_sr_v2_nrv_9_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_27_Im = FFT_sr_v2_nrv_9_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_28_Re = FFT_sr_v2_nrv_9_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_28_Im = FFT_sr_v2_nrv_9_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_29_Re = FFT_sr_v2_nrv_9_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_29_Im = FFT_sr_v2_nrv_9_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_30_Re = FFT_sr_v2_nrv_10_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_30_Im = FFT_sr_v2_nrv_10_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_31_Re = FFT_sr_v2_nrv_10_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_31_Im = FFT_sr_v2_nrv_10_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_32_Re = FFT_sr_v2_nrv_10_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_32_Im = FFT_sr_v2_nrv_10_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_33_Re = FFT_sr_v2_nrv_11_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_33_Im = FFT_sr_v2_nrv_11_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_34_Re = FFT_sr_v2_nrv_11_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_34_Im = FFT_sr_v2_nrv_11_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_35_Re = FFT_sr_v2_nrv_11_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_35_Im = FFT_sr_v2_nrv_11_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_36_Re = FFT_sr_v2_nrv_12_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_36_Im = FFT_sr_v2_nrv_12_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_37_Re = FFT_sr_v2_nrv_12_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_37_Im = FFT_sr_v2_nrv_12_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_38_Re = FFT_sr_v2_nrv_12_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_38_Im = FFT_sr_v2_nrv_12_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_39_Re = FFT_sr_v2_nrv_13_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_39_Im = FFT_sr_v2_nrv_13_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_40_Re = FFT_sr_v2_nrv_13_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_40_Im = FFT_sr_v2_nrv_13_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_41_Re = FFT_sr_v2_nrv_13_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_41_Im = FFT_sr_v2_nrv_13_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_42_Re = FFT_sr_v2_nrv_14_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_42_Im = FFT_sr_v2_nrv_14_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_43_Re = FFT_sr_v2_nrv_14_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_43_Im = FFT_sr_v2_nrv_14_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_44_Re = FFT_sr_v2_nrv_14_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_44_Im = FFT_sr_v2_nrv_14_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_45_Re = FFT_sr_v2_nrv_15_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_45_Im = FFT_sr_v2_nrv_15_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_46_Re = FFT_sr_v2_nrv_15_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_46_Im = FFT_sr_v2_nrv_15_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_47_Re = FFT_sr_v2_nrv_15_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_47_Im = FFT_sr_v2_nrv_15_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_48_Re = FFT_sr_v2_nrv_16_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_48_Im = FFT_sr_v2_nrv_16_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_49_Re = FFT_sr_v2_nrv_16_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_49_Im = FFT_sr_v2_nrv_16_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_50_Re = FFT_sr_v2_nrv_16_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_50_Im = FFT_sr_v2_nrv_16_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_51_Re = FFT_sr_v2_nrv_17_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_51_Im = FFT_sr_v2_nrv_17_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_52_Re = FFT_sr_v2_nrv_17_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_52_Im = FFT_sr_v2_nrv_17_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_53_Re = FFT_sr_v2_nrv_17_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_53_Im = FFT_sr_v2_nrv_17_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_54_Re = FFT_sr_v2_nrv_18_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_54_Im = FFT_sr_v2_nrv_18_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_55_Re = FFT_sr_v2_nrv_18_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_55_Im = FFT_sr_v2_nrv_18_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_56_Re = FFT_sr_v2_nrv_18_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_56_Im = FFT_sr_v2_nrv_18_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_57_Re = FFT_sr_v2_nrv_19_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_57_Im = FFT_sr_v2_nrv_19_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_58_Re = FFT_sr_v2_nrv_19_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_58_Im = FFT_sr_v2_nrv_19_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_59_Re = FFT_sr_v2_nrv_19_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_59_Im = FFT_sr_v2_nrv_19_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_60_Re = FFT_sr_v2_nrv_20_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_60_Im = FFT_sr_v2_nrv_20_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_61_Re = FFT_sr_v2_nrv_20_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_61_Im = FFT_sr_v2_nrv_20_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_62_Re = FFT_sr_v2_nrv_20_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_62_Im = FFT_sr_v2_nrv_20_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_63_Re = FFT_sr_v2_nrv_21_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_63_Im = FFT_sr_v2_nrv_21_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_64_Re = FFT_sr_v2_nrv_21_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_64_Im = FFT_sr_v2_nrv_21_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_65_Re = FFT_sr_v2_nrv_21_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_65_Im = FFT_sr_v2_nrv_21_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_66_Re = FFT_sr_v2_nrv_22_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_66_Im = FFT_sr_v2_nrv_22_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_67_Re = FFT_sr_v2_nrv_22_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_67_Im = FFT_sr_v2_nrv_22_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_68_Re = FFT_sr_v2_nrv_22_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_68_Im = FFT_sr_v2_nrv_22_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_69_Re = FFT_sr_v2_nrv_23_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_69_Im = FFT_sr_v2_nrv_23_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_70_Re = FFT_sr_v2_nrv_23_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_70_Im = FFT_sr_v2_nrv_23_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_71_Re = FFT_sr_v2_nrv_23_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_71_Im = FFT_sr_v2_nrv_23_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_72_Re = FFT_sr_v2_nrv_24_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_72_Im = FFT_sr_v2_nrv_24_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_73_Re = FFT_sr_v2_nrv_24_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_73_Im = FFT_sr_v2_nrv_24_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_74_Re = FFT_sr_v2_nrv_24_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_74_Im = FFT_sr_v2_nrv_24_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_75_Re = FFT_sr_v2_nrv_25_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_75_Im = FFT_sr_v2_nrv_25_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_76_Re = FFT_sr_v2_nrv_25_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_76_Im = FFT_sr_v2_nrv_25_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_77_Re = FFT_sr_v2_nrv_25_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_77_Im = FFT_sr_v2_nrv_25_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_78_Re = FFT_sr_v2_nrv_26_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_78_Im = FFT_sr_v2_nrv_26_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_79_Re = FFT_sr_v2_nrv_26_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_79_Im = FFT_sr_v2_nrv_26_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_80_Re = FFT_sr_v2_nrv_26_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_80_Im = FFT_sr_v2_nrv_26_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_81_Re = FFT_sr_v2_nrv_27_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_81_Im = FFT_sr_v2_nrv_27_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_82_Re = FFT_sr_v2_nrv_27_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_82_Im = FFT_sr_v2_nrv_27_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_83_Re = FFT_sr_v2_nrv_27_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_83_Im = FFT_sr_v2_nrv_27_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_84_Re = FFT_sr_v2_nrv_28_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_84_Im = FFT_sr_v2_nrv_28_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_85_Re = FFT_sr_v2_nrv_28_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_85_Im = FFT_sr_v2_nrv_28_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_86_Re = FFT_sr_v2_nrv_28_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_86_Im = FFT_sr_v2_nrv_28_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_87_Re = FFT_sr_v2_nrv_29_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_87_Im = FFT_sr_v2_nrv_29_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_88_Re = FFT_sr_v2_nrv_29_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_88_Im = FFT_sr_v2_nrv_29_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_89_Re = FFT_sr_v2_nrv_29_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_89_Im = FFT_sr_v2_nrv_29_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_90_Re = FFT_sr_v2_nrv_30_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_90_Im = FFT_sr_v2_nrv_30_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_91_Re = FFT_sr_v2_nrv_30_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_91_Im = FFT_sr_v2_nrv_30_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_92_Re = FFT_sr_v2_nrv_30_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_92_Im = FFT_sr_v2_nrv_30_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_93_Re = FFT_sr_v2_nrv_31_io_out_0_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_93_Im = FFT_sr_v2_nrv_31_io_out_0_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_94_Re = FFT_sr_v2_nrv_31_io_out_1_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_94_Im = FFT_sr_v2_nrv_31_io_out_1_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_95_Re = FFT_sr_v2_nrv_31_io_out_2_Re; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_1_io_in_95_Im = FFT_sr_v2_nrv_31_io_out_2_Im; // @[FFTDesigns.scala 3478:45]
  assign PermutationsBasic_2_io_in_0_Re = FFT_sr_v2_nrv_32_io_out_0_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_0_Im = FFT_sr_v2_nrv_32_io_out_0_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_1_Re = FFT_sr_v2_nrv_32_io_out_1_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_1_Im = FFT_sr_v2_nrv_32_io_out_1_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_2_Re = FFT_sr_v2_nrv_32_io_out_2_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_2_Im = FFT_sr_v2_nrv_32_io_out_2_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_3_Re = FFT_sr_v2_nrv_32_io_out_3_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_3_Im = FFT_sr_v2_nrv_32_io_out_3_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_4_Re = FFT_sr_v2_nrv_32_io_out_4_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_4_Im = FFT_sr_v2_nrv_32_io_out_4_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_5_Re = FFT_sr_v2_nrv_32_io_out_5_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_5_Im = FFT_sr_v2_nrv_32_io_out_5_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_6_Re = FFT_sr_v2_nrv_32_io_out_6_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_6_Im = FFT_sr_v2_nrv_32_io_out_6_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_7_Re = FFT_sr_v2_nrv_32_io_out_7_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_7_Im = FFT_sr_v2_nrv_32_io_out_7_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_8_Re = FFT_sr_v2_nrv_32_io_out_8_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_8_Im = FFT_sr_v2_nrv_32_io_out_8_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_9_Re = FFT_sr_v2_nrv_32_io_out_9_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_9_Im = FFT_sr_v2_nrv_32_io_out_9_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_10_Re = FFT_sr_v2_nrv_32_io_out_10_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_10_Im = FFT_sr_v2_nrv_32_io_out_10_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_11_Re = FFT_sr_v2_nrv_32_io_out_11_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_11_Im = FFT_sr_v2_nrv_32_io_out_11_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_12_Re = FFT_sr_v2_nrv_32_io_out_12_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_12_Im = FFT_sr_v2_nrv_32_io_out_12_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_13_Re = FFT_sr_v2_nrv_32_io_out_13_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_13_Im = FFT_sr_v2_nrv_32_io_out_13_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_14_Re = FFT_sr_v2_nrv_32_io_out_14_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_14_Im = FFT_sr_v2_nrv_32_io_out_14_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_15_Re = FFT_sr_v2_nrv_32_io_out_15_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_15_Im = FFT_sr_v2_nrv_32_io_out_15_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_16_Re = FFT_sr_v2_nrv_32_io_out_16_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_16_Im = FFT_sr_v2_nrv_32_io_out_16_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_17_Re = FFT_sr_v2_nrv_32_io_out_17_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_17_Im = FFT_sr_v2_nrv_32_io_out_17_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_18_Re = FFT_sr_v2_nrv_32_io_out_18_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_18_Im = FFT_sr_v2_nrv_32_io_out_18_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_19_Re = FFT_sr_v2_nrv_32_io_out_19_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_19_Im = FFT_sr_v2_nrv_32_io_out_19_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_20_Re = FFT_sr_v2_nrv_32_io_out_20_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_20_Im = FFT_sr_v2_nrv_32_io_out_20_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_21_Re = FFT_sr_v2_nrv_32_io_out_21_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_21_Im = FFT_sr_v2_nrv_32_io_out_21_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_22_Re = FFT_sr_v2_nrv_32_io_out_22_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_22_Im = FFT_sr_v2_nrv_32_io_out_22_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_23_Re = FFT_sr_v2_nrv_32_io_out_23_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_23_Im = FFT_sr_v2_nrv_32_io_out_23_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_24_Re = FFT_sr_v2_nrv_32_io_out_24_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_24_Im = FFT_sr_v2_nrv_32_io_out_24_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_25_Re = FFT_sr_v2_nrv_32_io_out_25_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_25_Im = FFT_sr_v2_nrv_32_io_out_25_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_26_Re = FFT_sr_v2_nrv_32_io_out_26_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_26_Im = FFT_sr_v2_nrv_32_io_out_26_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_27_Re = FFT_sr_v2_nrv_32_io_out_27_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_27_Im = FFT_sr_v2_nrv_32_io_out_27_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_28_Re = FFT_sr_v2_nrv_32_io_out_28_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_28_Im = FFT_sr_v2_nrv_32_io_out_28_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_29_Re = FFT_sr_v2_nrv_32_io_out_29_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_29_Im = FFT_sr_v2_nrv_32_io_out_29_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_30_Re = FFT_sr_v2_nrv_32_io_out_30_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_30_Im = FFT_sr_v2_nrv_32_io_out_30_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_31_Re = FFT_sr_v2_nrv_32_io_out_31_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_31_Im = FFT_sr_v2_nrv_32_io_out_31_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_32_Re = FFT_sr_v2_nrv_33_io_out_0_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_32_Im = FFT_sr_v2_nrv_33_io_out_0_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_33_Re = FFT_sr_v2_nrv_33_io_out_1_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_33_Im = FFT_sr_v2_nrv_33_io_out_1_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_34_Re = FFT_sr_v2_nrv_33_io_out_2_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_34_Im = FFT_sr_v2_nrv_33_io_out_2_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_35_Re = FFT_sr_v2_nrv_33_io_out_3_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_35_Im = FFT_sr_v2_nrv_33_io_out_3_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_36_Re = FFT_sr_v2_nrv_33_io_out_4_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_36_Im = FFT_sr_v2_nrv_33_io_out_4_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_37_Re = FFT_sr_v2_nrv_33_io_out_5_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_37_Im = FFT_sr_v2_nrv_33_io_out_5_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_38_Re = FFT_sr_v2_nrv_33_io_out_6_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_38_Im = FFT_sr_v2_nrv_33_io_out_6_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_39_Re = FFT_sr_v2_nrv_33_io_out_7_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_39_Im = FFT_sr_v2_nrv_33_io_out_7_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_40_Re = FFT_sr_v2_nrv_33_io_out_8_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_40_Im = FFT_sr_v2_nrv_33_io_out_8_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_41_Re = FFT_sr_v2_nrv_33_io_out_9_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_41_Im = FFT_sr_v2_nrv_33_io_out_9_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_42_Re = FFT_sr_v2_nrv_33_io_out_10_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_42_Im = FFT_sr_v2_nrv_33_io_out_10_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_43_Re = FFT_sr_v2_nrv_33_io_out_11_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_43_Im = FFT_sr_v2_nrv_33_io_out_11_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_44_Re = FFT_sr_v2_nrv_33_io_out_12_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_44_Im = FFT_sr_v2_nrv_33_io_out_12_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_45_Re = FFT_sr_v2_nrv_33_io_out_13_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_45_Im = FFT_sr_v2_nrv_33_io_out_13_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_46_Re = FFT_sr_v2_nrv_33_io_out_14_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_46_Im = FFT_sr_v2_nrv_33_io_out_14_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_47_Re = FFT_sr_v2_nrv_33_io_out_15_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_47_Im = FFT_sr_v2_nrv_33_io_out_15_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_48_Re = FFT_sr_v2_nrv_33_io_out_16_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_48_Im = FFT_sr_v2_nrv_33_io_out_16_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_49_Re = FFT_sr_v2_nrv_33_io_out_17_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_49_Im = FFT_sr_v2_nrv_33_io_out_17_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_50_Re = FFT_sr_v2_nrv_33_io_out_18_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_50_Im = FFT_sr_v2_nrv_33_io_out_18_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_51_Re = FFT_sr_v2_nrv_33_io_out_19_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_51_Im = FFT_sr_v2_nrv_33_io_out_19_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_52_Re = FFT_sr_v2_nrv_33_io_out_20_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_52_Im = FFT_sr_v2_nrv_33_io_out_20_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_53_Re = FFT_sr_v2_nrv_33_io_out_21_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_53_Im = FFT_sr_v2_nrv_33_io_out_21_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_54_Re = FFT_sr_v2_nrv_33_io_out_22_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_54_Im = FFT_sr_v2_nrv_33_io_out_22_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_55_Re = FFT_sr_v2_nrv_33_io_out_23_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_55_Im = FFT_sr_v2_nrv_33_io_out_23_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_56_Re = FFT_sr_v2_nrv_33_io_out_24_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_56_Im = FFT_sr_v2_nrv_33_io_out_24_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_57_Re = FFT_sr_v2_nrv_33_io_out_25_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_57_Im = FFT_sr_v2_nrv_33_io_out_25_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_58_Re = FFT_sr_v2_nrv_33_io_out_26_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_58_Im = FFT_sr_v2_nrv_33_io_out_26_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_59_Re = FFT_sr_v2_nrv_33_io_out_27_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_59_Im = FFT_sr_v2_nrv_33_io_out_27_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_60_Re = FFT_sr_v2_nrv_33_io_out_28_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_60_Im = FFT_sr_v2_nrv_33_io_out_28_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_61_Re = FFT_sr_v2_nrv_33_io_out_29_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_61_Im = FFT_sr_v2_nrv_33_io_out_29_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_62_Re = FFT_sr_v2_nrv_33_io_out_30_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_62_Im = FFT_sr_v2_nrv_33_io_out_30_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_63_Re = FFT_sr_v2_nrv_33_io_out_31_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_63_Im = FFT_sr_v2_nrv_33_io_out_31_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_64_Re = FFT_sr_v2_nrv_34_io_out_0_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_64_Im = FFT_sr_v2_nrv_34_io_out_0_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_65_Re = FFT_sr_v2_nrv_34_io_out_1_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_65_Im = FFT_sr_v2_nrv_34_io_out_1_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_66_Re = FFT_sr_v2_nrv_34_io_out_2_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_66_Im = FFT_sr_v2_nrv_34_io_out_2_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_67_Re = FFT_sr_v2_nrv_34_io_out_3_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_67_Im = FFT_sr_v2_nrv_34_io_out_3_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_68_Re = FFT_sr_v2_nrv_34_io_out_4_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_68_Im = FFT_sr_v2_nrv_34_io_out_4_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_69_Re = FFT_sr_v2_nrv_34_io_out_5_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_69_Im = FFT_sr_v2_nrv_34_io_out_5_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_70_Re = FFT_sr_v2_nrv_34_io_out_6_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_70_Im = FFT_sr_v2_nrv_34_io_out_6_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_71_Re = FFT_sr_v2_nrv_34_io_out_7_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_71_Im = FFT_sr_v2_nrv_34_io_out_7_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_72_Re = FFT_sr_v2_nrv_34_io_out_8_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_72_Im = FFT_sr_v2_nrv_34_io_out_8_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_73_Re = FFT_sr_v2_nrv_34_io_out_9_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_73_Im = FFT_sr_v2_nrv_34_io_out_9_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_74_Re = FFT_sr_v2_nrv_34_io_out_10_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_74_Im = FFT_sr_v2_nrv_34_io_out_10_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_75_Re = FFT_sr_v2_nrv_34_io_out_11_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_75_Im = FFT_sr_v2_nrv_34_io_out_11_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_76_Re = FFT_sr_v2_nrv_34_io_out_12_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_76_Im = FFT_sr_v2_nrv_34_io_out_12_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_77_Re = FFT_sr_v2_nrv_34_io_out_13_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_77_Im = FFT_sr_v2_nrv_34_io_out_13_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_78_Re = FFT_sr_v2_nrv_34_io_out_14_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_78_Im = FFT_sr_v2_nrv_34_io_out_14_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_79_Re = FFT_sr_v2_nrv_34_io_out_15_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_79_Im = FFT_sr_v2_nrv_34_io_out_15_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_80_Re = FFT_sr_v2_nrv_34_io_out_16_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_80_Im = FFT_sr_v2_nrv_34_io_out_16_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_81_Re = FFT_sr_v2_nrv_34_io_out_17_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_81_Im = FFT_sr_v2_nrv_34_io_out_17_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_82_Re = FFT_sr_v2_nrv_34_io_out_18_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_82_Im = FFT_sr_v2_nrv_34_io_out_18_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_83_Re = FFT_sr_v2_nrv_34_io_out_19_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_83_Im = FFT_sr_v2_nrv_34_io_out_19_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_84_Re = FFT_sr_v2_nrv_34_io_out_20_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_84_Im = FFT_sr_v2_nrv_34_io_out_20_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_85_Re = FFT_sr_v2_nrv_34_io_out_21_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_85_Im = FFT_sr_v2_nrv_34_io_out_21_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_86_Re = FFT_sr_v2_nrv_34_io_out_22_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_86_Im = FFT_sr_v2_nrv_34_io_out_22_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_87_Re = FFT_sr_v2_nrv_34_io_out_23_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_87_Im = FFT_sr_v2_nrv_34_io_out_23_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_88_Re = FFT_sr_v2_nrv_34_io_out_24_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_88_Im = FFT_sr_v2_nrv_34_io_out_24_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_89_Re = FFT_sr_v2_nrv_34_io_out_25_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_89_Im = FFT_sr_v2_nrv_34_io_out_25_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_90_Re = FFT_sr_v2_nrv_34_io_out_26_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_90_Im = FFT_sr_v2_nrv_34_io_out_26_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_91_Re = FFT_sr_v2_nrv_34_io_out_27_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_91_Im = FFT_sr_v2_nrv_34_io_out_27_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_92_Re = FFT_sr_v2_nrv_34_io_out_28_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_92_Im = FFT_sr_v2_nrv_34_io_out_28_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_93_Re = FFT_sr_v2_nrv_34_io_out_29_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_93_Im = FFT_sr_v2_nrv_34_io_out_29_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_94_Re = FFT_sr_v2_nrv_34_io_out_30_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_94_Im = FFT_sr_v2_nrv_34_io_out_30_Im; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_95_Re = FFT_sr_v2_nrv_34_io_out_31_Re; // @[FFTDesigns.scala 3480:45]
  assign PermutationsBasic_2_io_in_95_Im = FFT_sr_v2_nrv_34_io_out_31_Im; // @[FFTDesigns.scala 3480:45]
  assign TwiddleFactors_mr_clock = clock;
  assign TwiddleFactors_mr_reset = reset;
  assign TwiddleFactors_mr_io_in_0_Re = PermutationsBasic_1_io_out_0_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_0_Im = PermutationsBasic_1_io_out_0_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_1_Re = PermutationsBasic_1_io_out_1_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_1_Im = PermutationsBasic_1_io_out_1_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_2_Re = PermutationsBasic_1_io_out_2_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_2_Im = PermutationsBasic_1_io_out_2_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_3_Re = PermutationsBasic_1_io_out_3_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_3_Im = PermutationsBasic_1_io_out_3_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_4_Re = PermutationsBasic_1_io_out_4_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_4_Im = PermutationsBasic_1_io_out_4_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_5_Re = PermutationsBasic_1_io_out_5_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_5_Im = PermutationsBasic_1_io_out_5_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_6_Re = PermutationsBasic_1_io_out_6_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_6_Im = PermutationsBasic_1_io_out_6_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_7_Re = PermutationsBasic_1_io_out_7_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_7_Im = PermutationsBasic_1_io_out_7_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_8_Re = PermutationsBasic_1_io_out_8_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_8_Im = PermutationsBasic_1_io_out_8_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_9_Re = PermutationsBasic_1_io_out_9_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_9_Im = PermutationsBasic_1_io_out_9_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_10_Re = PermutationsBasic_1_io_out_10_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_10_Im = PermutationsBasic_1_io_out_10_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_11_Re = PermutationsBasic_1_io_out_11_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_11_Im = PermutationsBasic_1_io_out_11_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_12_Re = PermutationsBasic_1_io_out_12_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_12_Im = PermutationsBasic_1_io_out_12_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_13_Re = PermutationsBasic_1_io_out_13_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_13_Im = PermutationsBasic_1_io_out_13_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_14_Re = PermutationsBasic_1_io_out_14_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_14_Im = PermutationsBasic_1_io_out_14_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_15_Re = PermutationsBasic_1_io_out_15_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_15_Im = PermutationsBasic_1_io_out_15_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_16_Re = PermutationsBasic_1_io_out_16_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_16_Im = PermutationsBasic_1_io_out_16_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_17_Re = PermutationsBasic_1_io_out_17_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_17_Im = PermutationsBasic_1_io_out_17_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_18_Re = PermutationsBasic_1_io_out_18_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_18_Im = PermutationsBasic_1_io_out_18_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_19_Re = PermutationsBasic_1_io_out_19_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_19_Im = PermutationsBasic_1_io_out_19_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_20_Re = PermutationsBasic_1_io_out_20_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_20_Im = PermutationsBasic_1_io_out_20_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_21_Re = PermutationsBasic_1_io_out_21_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_21_Im = PermutationsBasic_1_io_out_21_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_22_Re = PermutationsBasic_1_io_out_22_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_22_Im = PermutationsBasic_1_io_out_22_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_23_Re = PermutationsBasic_1_io_out_23_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_23_Im = PermutationsBasic_1_io_out_23_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_24_Re = PermutationsBasic_1_io_out_24_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_24_Im = PermutationsBasic_1_io_out_24_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_25_Re = PermutationsBasic_1_io_out_25_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_25_Im = PermutationsBasic_1_io_out_25_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_26_Re = PermutationsBasic_1_io_out_26_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_26_Im = PermutationsBasic_1_io_out_26_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_27_Re = PermutationsBasic_1_io_out_27_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_27_Im = PermutationsBasic_1_io_out_27_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_28_Re = PermutationsBasic_1_io_out_28_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_28_Im = PermutationsBasic_1_io_out_28_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_29_Re = PermutationsBasic_1_io_out_29_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_29_Im = PermutationsBasic_1_io_out_29_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_30_Re = PermutationsBasic_1_io_out_30_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_30_Im = PermutationsBasic_1_io_out_30_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_31_Re = PermutationsBasic_1_io_out_31_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_31_Im = PermutationsBasic_1_io_out_31_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_32_Re = PermutationsBasic_1_io_out_32_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_32_Im = PermutationsBasic_1_io_out_32_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_33_Re = PermutationsBasic_1_io_out_33_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_33_Im = PermutationsBasic_1_io_out_33_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_34_Re = PermutationsBasic_1_io_out_34_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_34_Im = PermutationsBasic_1_io_out_34_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_35_Re = PermutationsBasic_1_io_out_35_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_35_Im = PermutationsBasic_1_io_out_35_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_36_Re = PermutationsBasic_1_io_out_36_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_36_Im = PermutationsBasic_1_io_out_36_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_37_Re = PermutationsBasic_1_io_out_37_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_37_Im = PermutationsBasic_1_io_out_37_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_38_Re = PermutationsBasic_1_io_out_38_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_38_Im = PermutationsBasic_1_io_out_38_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_39_Re = PermutationsBasic_1_io_out_39_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_39_Im = PermutationsBasic_1_io_out_39_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_40_Re = PermutationsBasic_1_io_out_40_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_40_Im = PermutationsBasic_1_io_out_40_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_41_Re = PermutationsBasic_1_io_out_41_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_41_Im = PermutationsBasic_1_io_out_41_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_42_Re = PermutationsBasic_1_io_out_42_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_42_Im = PermutationsBasic_1_io_out_42_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_43_Re = PermutationsBasic_1_io_out_43_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_43_Im = PermutationsBasic_1_io_out_43_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_44_Re = PermutationsBasic_1_io_out_44_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_44_Im = PermutationsBasic_1_io_out_44_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_45_Re = PermutationsBasic_1_io_out_45_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_45_Im = PermutationsBasic_1_io_out_45_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_46_Re = PermutationsBasic_1_io_out_46_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_46_Im = PermutationsBasic_1_io_out_46_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_47_Re = PermutationsBasic_1_io_out_47_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_47_Im = PermutationsBasic_1_io_out_47_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_48_Re = PermutationsBasic_1_io_out_48_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_48_Im = PermutationsBasic_1_io_out_48_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_49_Re = PermutationsBasic_1_io_out_49_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_49_Im = PermutationsBasic_1_io_out_49_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_50_Re = PermutationsBasic_1_io_out_50_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_50_Im = PermutationsBasic_1_io_out_50_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_51_Re = PermutationsBasic_1_io_out_51_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_51_Im = PermutationsBasic_1_io_out_51_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_52_Re = PermutationsBasic_1_io_out_52_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_52_Im = PermutationsBasic_1_io_out_52_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_53_Re = PermutationsBasic_1_io_out_53_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_53_Im = PermutationsBasic_1_io_out_53_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_54_Re = PermutationsBasic_1_io_out_54_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_54_Im = PermutationsBasic_1_io_out_54_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_55_Re = PermutationsBasic_1_io_out_55_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_55_Im = PermutationsBasic_1_io_out_55_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_56_Re = PermutationsBasic_1_io_out_56_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_56_Im = PermutationsBasic_1_io_out_56_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_57_Re = PermutationsBasic_1_io_out_57_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_57_Im = PermutationsBasic_1_io_out_57_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_58_Re = PermutationsBasic_1_io_out_58_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_58_Im = PermutationsBasic_1_io_out_58_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_59_Re = PermutationsBasic_1_io_out_59_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_59_Im = PermutationsBasic_1_io_out_59_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_60_Re = PermutationsBasic_1_io_out_60_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_60_Im = PermutationsBasic_1_io_out_60_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_61_Re = PermutationsBasic_1_io_out_61_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_61_Im = PermutationsBasic_1_io_out_61_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_62_Re = PermutationsBasic_1_io_out_62_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_62_Im = PermutationsBasic_1_io_out_62_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_63_Re = PermutationsBasic_1_io_out_63_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_63_Im = PermutationsBasic_1_io_out_63_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_64_Re = PermutationsBasic_1_io_out_64_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_64_Im = PermutationsBasic_1_io_out_64_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_65_Re = PermutationsBasic_1_io_out_65_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_65_Im = PermutationsBasic_1_io_out_65_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_66_Re = PermutationsBasic_1_io_out_66_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_66_Im = PermutationsBasic_1_io_out_66_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_67_Re = PermutationsBasic_1_io_out_67_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_67_Im = PermutationsBasic_1_io_out_67_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_68_Re = PermutationsBasic_1_io_out_68_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_68_Im = PermutationsBasic_1_io_out_68_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_69_Re = PermutationsBasic_1_io_out_69_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_69_Im = PermutationsBasic_1_io_out_69_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_70_Re = PermutationsBasic_1_io_out_70_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_70_Im = PermutationsBasic_1_io_out_70_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_71_Re = PermutationsBasic_1_io_out_71_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_71_Im = PermutationsBasic_1_io_out_71_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_72_Re = PermutationsBasic_1_io_out_72_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_72_Im = PermutationsBasic_1_io_out_72_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_73_Re = PermutationsBasic_1_io_out_73_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_73_Im = PermutationsBasic_1_io_out_73_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_74_Re = PermutationsBasic_1_io_out_74_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_74_Im = PermutationsBasic_1_io_out_74_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_75_Re = PermutationsBasic_1_io_out_75_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_75_Im = PermutationsBasic_1_io_out_75_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_76_Re = PermutationsBasic_1_io_out_76_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_76_Im = PermutationsBasic_1_io_out_76_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_77_Re = PermutationsBasic_1_io_out_77_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_77_Im = PermutationsBasic_1_io_out_77_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_78_Re = PermutationsBasic_1_io_out_78_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_78_Im = PermutationsBasic_1_io_out_78_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_79_Re = PermutationsBasic_1_io_out_79_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_79_Im = PermutationsBasic_1_io_out_79_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_80_Re = PermutationsBasic_1_io_out_80_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_80_Im = PermutationsBasic_1_io_out_80_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_81_Re = PermutationsBasic_1_io_out_81_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_81_Im = PermutationsBasic_1_io_out_81_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_82_Re = PermutationsBasic_1_io_out_82_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_82_Im = PermutationsBasic_1_io_out_82_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_83_Re = PermutationsBasic_1_io_out_83_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_83_Im = PermutationsBasic_1_io_out_83_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_84_Re = PermutationsBasic_1_io_out_84_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_84_Im = PermutationsBasic_1_io_out_84_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_85_Re = PermutationsBasic_1_io_out_85_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_85_Im = PermutationsBasic_1_io_out_85_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_86_Re = PermutationsBasic_1_io_out_86_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_86_Im = PermutationsBasic_1_io_out_86_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_87_Re = PermutationsBasic_1_io_out_87_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_87_Im = PermutationsBasic_1_io_out_87_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_88_Re = PermutationsBasic_1_io_out_88_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_88_Im = PermutationsBasic_1_io_out_88_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_89_Re = PermutationsBasic_1_io_out_89_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_89_Im = PermutationsBasic_1_io_out_89_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_90_Re = PermutationsBasic_1_io_out_90_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_90_Im = PermutationsBasic_1_io_out_90_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_91_Re = PermutationsBasic_1_io_out_91_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_91_Im = PermutationsBasic_1_io_out_91_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_92_Re = PermutationsBasic_1_io_out_92_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_92_Im = PermutationsBasic_1_io_out_92_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_93_Re = PermutationsBasic_1_io_out_93_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_93_Im = PermutationsBasic_1_io_out_93_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_94_Re = PermutationsBasic_1_io_out_94_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_94_Im = PermutationsBasic_1_io_out_94_Im; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_95_Re = PermutationsBasic_1_io_out_95_Re; // @[FFTDesigns.scala 3462:20]
  assign TwiddleFactors_mr_io_in_95_Im = PermutationsBasic_1_io_out_95_Im; // @[FFTDesigns.scala 3462:20]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_0 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_0 <= io_in_ready; // @[FFTDesigns.scala 3430:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_1 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_1 <= regdelays_0; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_2 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_2 <= regdelays_1; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_3 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_3 <= regdelays_2; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_4 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_4 <= regdelays_3; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_5 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_5 <= regdelays_4; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_6 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_6 <= regdelays_5; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_7 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_7 <= regdelays_6; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_8 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_8 <= regdelays_7; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_9 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_9 <= regdelays_8; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_10 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_10 <= regdelays_9; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_11 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_11 <= regdelays_10; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_12 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_12 <= regdelays_11; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_13 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_13 <= regdelays_12; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_14 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_14 <= regdelays_13; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_15 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_15 <= regdelays_14; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3427:28]
      regdelays_16 <= 1'h0; // @[FFTDesigns.scala 3427:28]
    end else begin
      regdelays_16 <= regdelays_15; // @[FFTDesigns.scala 3432:22]
    end
    if (reset) begin // @[FFTDesigns.scala 3435:31]
      out_regdelay <= 1'h0; // @[FFTDesigns.scala 3435:31]
    end else begin
      out_regdelay <= regdelays_16;
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_0_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_0_Re <= PermutationsBasic_2_io_out_0_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_0_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_0_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_0_Im <= PermutationsBasic_2_io_out_0_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_0_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_1_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_1_Re <= PermutationsBasic_2_io_out_1_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_1_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_1_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_1_Im <= PermutationsBasic_2_io_out_1_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_1_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_2_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_2_Re <= PermutationsBasic_2_io_out_2_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_2_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_2_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_2_Im <= PermutationsBasic_2_io_out_2_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_2_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_3_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_3_Re <= PermutationsBasic_2_io_out_3_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_3_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_3_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_3_Im <= PermutationsBasic_2_io_out_3_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_3_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_4_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_4_Re <= PermutationsBasic_2_io_out_4_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_4_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_4_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_4_Im <= PermutationsBasic_2_io_out_4_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_4_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_5_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_5_Re <= PermutationsBasic_2_io_out_5_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_5_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_5_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_5_Im <= PermutationsBasic_2_io_out_5_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_5_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_6_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_6_Re <= PermutationsBasic_2_io_out_6_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_6_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_6_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_6_Im <= PermutationsBasic_2_io_out_6_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_6_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_7_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_7_Re <= PermutationsBasic_2_io_out_7_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_7_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_7_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_7_Im <= PermutationsBasic_2_io_out_7_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_7_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_8_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_8_Re <= PermutationsBasic_2_io_out_8_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_8_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_8_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_8_Im <= PermutationsBasic_2_io_out_8_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_8_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_9_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_9_Re <= PermutationsBasic_2_io_out_9_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_9_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_9_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_9_Im <= PermutationsBasic_2_io_out_9_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_9_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_10_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_10_Re <= PermutationsBasic_2_io_out_10_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_10_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_10_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_10_Im <= PermutationsBasic_2_io_out_10_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_10_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_11_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_11_Re <= PermutationsBasic_2_io_out_11_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_11_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_11_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_11_Im <= PermutationsBasic_2_io_out_11_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_11_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_12_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_12_Re <= PermutationsBasic_2_io_out_12_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_12_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_12_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_12_Im <= PermutationsBasic_2_io_out_12_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_12_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_13_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_13_Re <= PermutationsBasic_2_io_out_13_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_13_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_13_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_13_Im <= PermutationsBasic_2_io_out_13_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_13_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_14_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_14_Re <= PermutationsBasic_2_io_out_14_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_14_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_14_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_14_Im <= PermutationsBasic_2_io_out_14_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_14_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_15_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_15_Re <= PermutationsBasic_2_io_out_15_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_15_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_15_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_15_Im <= PermutationsBasic_2_io_out_15_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_15_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_16_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_16_Re <= PermutationsBasic_2_io_out_16_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_16_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_16_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_16_Im <= PermutationsBasic_2_io_out_16_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_16_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_17_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_17_Re <= PermutationsBasic_2_io_out_17_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_17_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_17_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_17_Im <= PermutationsBasic_2_io_out_17_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_17_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_18_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_18_Re <= PermutationsBasic_2_io_out_18_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_18_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_18_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_18_Im <= PermutationsBasic_2_io_out_18_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_18_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_19_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_19_Re <= PermutationsBasic_2_io_out_19_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_19_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_19_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_19_Im <= PermutationsBasic_2_io_out_19_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_19_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_20_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_20_Re <= PermutationsBasic_2_io_out_20_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_20_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_20_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_20_Im <= PermutationsBasic_2_io_out_20_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_20_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_21_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_21_Re <= PermutationsBasic_2_io_out_21_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_21_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_21_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_21_Im <= PermutationsBasic_2_io_out_21_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_21_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_22_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_22_Re <= PermutationsBasic_2_io_out_22_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_22_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_22_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_22_Im <= PermutationsBasic_2_io_out_22_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_22_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_23_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_23_Re <= PermutationsBasic_2_io_out_23_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_23_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_23_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_23_Im <= PermutationsBasic_2_io_out_23_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_23_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_24_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_24_Re <= PermutationsBasic_2_io_out_24_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_24_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_24_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_24_Im <= PermutationsBasic_2_io_out_24_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_24_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_25_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_25_Re <= PermutationsBasic_2_io_out_25_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_25_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_25_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_25_Im <= PermutationsBasic_2_io_out_25_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_25_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_26_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_26_Re <= PermutationsBasic_2_io_out_26_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_26_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_26_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_26_Im <= PermutationsBasic_2_io_out_26_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_26_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_27_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_27_Re <= PermutationsBasic_2_io_out_27_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_27_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_27_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_27_Im <= PermutationsBasic_2_io_out_27_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_27_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_28_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_28_Re <= PermutationsBasic_2_io_out_28_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_28_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_28_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_28_Im <= PermutationsBasic_2_io_out_28_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_28_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_29_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_29_Re <= PermutationsBasic_2_io_out_29_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_29_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_29_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_29_Im <= PermutationsBasic_2_io_out_29_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_29_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_30_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_30_Re <= PermutationsBasic_2_io_out_30_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_30_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_30_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_30_Im <= PermutationsBasic_2_io_out_30_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_30_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_31_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_31_Re <= PermutationsBasic_2_io_out_31_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_31_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_31_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_31_Im <= PermutationsBasic_2_io_out_31_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_31_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_32_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_32_Re <= PermutationsBasic_2_io_out_32_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_32_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_32_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_32_Im <= PermutationsBasic_2_io_out_32_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_32_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_33_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_33_Re <= PermutationsBasic_2_io_out_33_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_33_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_33_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_33_Im <= PermutationsBasic_2_io_out_33_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_33_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_34_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_34_Re <= PermutationsBasic_2_io_out_34_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_34_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_34_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_34_Im <= PermutationsBasic_2_io_out_34_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_34_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_35_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_35_Re <= PermutationsBasic_2_io_out_35_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_35_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_35_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_35_Im <= PermutationsBasic_2_io_out_35_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_35_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_36_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_36_Re <= PermutationsBasic_2_io_out_36_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_36_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_36_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_36_Im <= PermutationsBasic_2_io_out_36_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_36_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_37_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_37_Re <= PermutationsBasic_2_io_out_37_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_37_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_37_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_37_Im <= PermutationsBasic_2_io_out_37_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_37_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_38_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_38_Re <= PermutationsBasic_2_io_out_38_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_38_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_38_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_38_Im <= PermutationsBasic_2_io_out_38_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_38_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_39_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_39_Re <= PermutationsBasic_2_io_out_39_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_39_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_39_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_39_Im <= PermutationsBasic_2_io_out_39_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_39_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_40_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_40_Re <= PermutationsBasic_2_io_out_40_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_40_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_40_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_40_Im <= PermutationsBasic_2_io_out_40_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_40_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_41_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_41_Re <= PermutationsBasic_2_io_out_41_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_41_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_41_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_41_Im <= PermutationsBasic_2_io_out_41_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_41_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_42_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_42_Re <= PermutationsBasic_2_io_out_42_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_42_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_42_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_42_Im <= PermutationsBasic_2_io_out_42_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_42_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_43_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_43_Re <= PermutationsBasic_2_io_out_43_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_43_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_43_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_43_Im <= PermutationsBasic_2_io_out_43_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_43_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_44_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_44_Re <= PermutationsBasic_2_io_out_44_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_44_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_44_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_44_Im <= PermutationsBasic_2_io_out_44_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_44_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_45_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_45_Re <= PermutationsBasic_2_io_out_45_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_45_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_45_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_45_Im <= PermutationsBasic_2_io_out_45_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_45_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_46_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_46_Re <= PermutationsBasic_2_io_out_46_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_46_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_46_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_46_Im <= PermutationsBasic_2_io_out_46_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_46_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_47_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_47_Re <= PermutationsBasic_2_io_out_47_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_47_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_47_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_47_Im <= PermutationsBasic_2_io_out_47_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_47_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_48_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_48_Re <= PermutationsBasic_2_io_out_48_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_48_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_48_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_48_Im <= PermutationsBasic_2_io_out_48_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_48_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_49_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_49_Re <= PermutationsBasic_2_io_out_49_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_49_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_49_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_49_Im <= PermutationsBasic_2_io_out_49_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_49_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_50_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_50_Re <= PermutationsBasic_2_io_out_50_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_50_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_50_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_50_Im <= PermutationsBasic_2_io_out_50_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_50_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_51_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_51_Re <= PermutationsBasic_2_io_out_51_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_51_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_51_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_51_Im <= PermutationsBasic_2_io_out_51_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_51_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_52_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_52_Re <= PermutationsBasic_2_io_out_52_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_52_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_52_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_52_Im <= PermutationsBasic_2_io_out_52_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_52_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_53_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_53_Re <= PermutationsBasic_2_io_out_53_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_53_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_53_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_53_Im <= PermutationsBasic_2_io_out_53_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_53_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_54_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_54_Re <= PermutationsBasic_2_io_out_54_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_54_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_54_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_54_Im <= PermutationsBasic_2_io_out_54_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_54_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_55_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_55_Re <= PermutationsBasic_2_io_out_55_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_55_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_55_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_55_Im <= PermutationsBasic_2_io_out_55_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_55_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_56_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_56_Re <= PermutationsBasic_2_io_out_56_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_56_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_56_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_56_Im <= PermutationsBasic_2_io_out_56_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_56_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_57_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_57_Re <= PermutationsBasic_2_io_out_57_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_57_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_57_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_57_Im <= PermutationsBasic_2_io_out_57_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_57_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_58_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_58_Re <= PermutationsBasic_2_io_out_58_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_58_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_58_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_58_Im <= PermutationsBasic_2_io_out_58_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_58_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_59_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_59_Re <= PermutationsBasic_2_io_out_59_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_59_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_59_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_59_Im <= PermutationsBasic_2_io_out_59_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_59_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_60_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_60_Re <= PermutationsBasic_2_io_out_60_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_60_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_60_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_60_Im <= PermutationsBasic_2_io_out_60_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_60_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_61_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_61_Re <= PermutationsBasic_2_io_out_61_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_61_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_61_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_61_Im <= PermutationsBasic_2_io_out_61_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_61_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_62_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_62_Re <= PermutationsBasic_2_io_out_62_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_62_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_62_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_62_Im <= PermutationsBasic_2_io_out_62_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_62_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_63_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_63_Re <= PermutationsBasic_2_io_out_63_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_63_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_63_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_63_Im <= PermutationsBasic_2_io_out_63_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_63_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_64_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_64_Re <= PermutationsBasic_2_io_out_64_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_64_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_64_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_64_Im <= PermutationsBasic_2_io_out_64_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_64_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_65_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_65_Re <= PermutationsBasic_2_io_out_65_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_65_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_65_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_65_Im <= PermutationsBasic_2_io_out_65_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_65_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_66_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_66_Re <= PermutationsBasic_2_io_out_66_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_66_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_66_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_66_Im <= PermutationsBasic_2_io_out_66_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_66_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_67_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_67_Re <= PermutationsBasic_2_io_out_67_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_67_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_67_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_67_Im <= PermutationsBasic_2_io_out_67_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_67_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_68_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_68_Re <= PermutationsBasic_2_io_out_68_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_68_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_68_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_68_Im <= PermutationsBasic_2_io_out_68_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_68_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_69_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_69_Re <= PermutationsBasic_2_io_out_69_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_69_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_69_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_69_Im <= PermutationsBasic_2_io_out_69_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_69_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_70_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_70_Re <= PermutationsBasic_2_io_out_70_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_70_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_70_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_70_Im <= PermutationsBasic_2_io_out_70_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_70_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_71_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_71_Re <= PermutationsBasic_2_io_out_71_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_71_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_71_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_71_Im <= PermutationsBasic_2_io_out_71_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_71_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_72_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_72_Re <= PermutationsBasic_2_io_out_72_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_72_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_72_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_72_Im <= PermutationsBasic_2_io_out_72_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_72_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_73_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_73_Re <= PermutationsBasic_2_io_out_73_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_73_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_73_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_73_Im <= PermutationsBasic_2_io_out_73_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_73_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_74_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_74_Re <= PermutationsBasic_2_io_out_74_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_74_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_74_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_74_Im <= PermutationsBasic_2_io_out_74_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_74_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_75_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_75_Re <= PermutationsBasic_2_io_out_75_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_75_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_75_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_75_Im <= PermutationsBasic_2_io_out_75_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_75_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_76_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_76_Re <= PermutationsBasic_2_io_out_76_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_76_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_76_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_76_Im <= PermutationsBasic_2_io_out_76_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_76_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_77_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_77_Re <= PermutationsBasic_2_io_out_77_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_77_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_77_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_77_Im <= PermutationsBasic_2_io_out_77_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_77_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_78_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_78_Re <= PermutationsBasic_2_io_out_78_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_78_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_78_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_78_Im <= PermutationsBasic_2_io_out_78_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_78_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_79_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_79_Re <= PermutationsBasic_2_io_out_79_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_79_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_79_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_79_Im <= PermutationsBasic_2_io_out_79_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_79_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_80_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_80_Re <= PermutationsBasic_2_io_out_80_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_80_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_80_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_80_Im <= PermutationsBasic_2_io_out_80_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_80_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_81_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_81_Re <= PermutationsBasic_2_io_out_81_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_81_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_81_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_81_Im <= PermutationsBasic_2_io_out_81_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_81_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_82_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_82_Re <= PermutationsBasic_2_io_out_82_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_82_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_82_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_82_Im <= PermutationsBasic_2_io_out_82_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_82_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_83_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_83_Re <= PermutationsBasic_2_io_out_83_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_83_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_83_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_83_Im <= PermutationsBasic_2_io_out_83_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_83_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_84_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_84_Re <= PermutationsBasic_2_io_out_84_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_84_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_84_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_84_Im <= PermutationsBasic_2_io_out_84_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_84_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_85_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_85_Re <= PermutationsBasic_2_io_out_85_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_85_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_85_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_85_Im <= PermutationsBasic_2_io_out_85_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_85_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_86_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_86_Re <= PermutationsBasic_2_io_out_86_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_86_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_86_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_86_Im <= PermutationsBasic_2_io_out_86_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_86_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_87_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_87_Re <= PermutationsBasic_2_io_out_87_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_87_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_87_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_87_Im <= PermutationsBasic_2_io_out_87_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_87_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_88_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_88_Re <= PermutationsBasic_2_io_out_88_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_88_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_88_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_88_Im <= PermutationsBasic_2_io_out_88_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_88_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_89_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_89_Re <= PermutationsBasic_2_io_out_89_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_89_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_89_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_89_Im <= PermutationsBasic_2_io_out_89_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_89_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_90_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_90_Re <= PermutationsBasic_2_io_out_90_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_90_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_90_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_90_Im <= PermutationsBasic_2_io_out_90_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_90_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_91_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_91_Re <= PermutationsBasic_2_io_out_91_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_91_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_91_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_91_Im <= PermutationsBasic_2_io_out_91_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_91_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_92_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_92_Re <= PermutationsBasic_2_io_out_92_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_92_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_92_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_92_Im <= PermutationsBasic_2_io_out_92_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_92_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_93_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_93_Re <= PermutationsBasic_2_io_out_93_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_93_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_93_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_93_Im <= PermutationsBasic_2_io_out_93_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_93_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_94_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_94_Re <= PermutationsBasic_2_io_out_94_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_94_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_94_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_94_Im <= PermutationsBasic_2_io_out_94_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_94_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_95_Re <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_95_Re <= PermutationsBasic_2_io_out_95_Re; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_95_Re <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
    if (reset) begin // @[FFTDesigns.scala 3463:30]
      out_results_95_Im <= 32'h0; // @[FFTDesigns.scala 3463:30]
    end else if (regdelays_16) begin // @[FFTDesigns.scala 3464:37]
      out_results_95_Im <= PermutationsBasic_2_io_out_95_Im; // @[FFTDesigns.scala 3465:19]
    end else begin
      out_results_95_Im <= 32'h0; // @[FFTDesigns.scala 3469:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regdelays_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  regdelays_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  regdelays_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  regdelays_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  regdelays_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  regdelays_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  regdelays_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  regdelays_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  regdelays_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  regdelays_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  regdelays_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  regdelays_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  regdelays_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  regdelays_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  regdelays_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  regdelays_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  regdelays_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  out_regdelay = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  out_results_0_Re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  out_results_0_Im = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  out_results_1_Re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  out_results_1_Im = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  out_results_2_Re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  out_results_2_Im = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  out_results_3_Re = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  out_results_3_Im = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  out_results_4_Re = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  out_results_4_Im = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  out_results_5_Re = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  out_results_5_Im = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  out_results_6_Re = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  out_results_6_Im = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  out_results_7_Re = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  out_results_7_Im = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  out_results_8_Re = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  out_results_8_Im = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  out_results_9_Re = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  out_results_9_Im = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  out_results_10_Re = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  out_results_10_Im = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  out_results_11_Re = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  out_results_11_Im = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  out_results_12_Re = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  out_results_12_Im = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  out_results_13_Re = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  out_results_13_Im = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  out_results_14_Re = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  out_results_14_Im = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  out_results_15_Re = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  out_results_15_Im = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  out_results_16_Re = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  out_results_16_Im = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  out_results_17_Re = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  out_results_17_Im = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  out_results_18_Re = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  out_results_18_Im = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  out_results_19_Re = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  out_results_19_Im = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  out_results_20_Re = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  out_results_20_Im = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  out_results_21_Re = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  out_results_21_Im = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  out_results_22_Re = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  out_results_22_Im = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  out_results_23_Re = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  out_results_23_Im = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  out_results_24_Re = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  out_results_24_Im = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  out_results_25_Re = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  out_results_25_Im = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  out_results_26_Re = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  out_results_26_Im = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  out_results_27_Re = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  out_results_27_Im = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  out_results_28_Re = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  out_results_28_Im = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  out_results_29_Re = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  out_results_29_Im = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  out_results_30_Re = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  out_results_30_Im = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  out_results_31_Re = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  out_results_31_Im = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  out_results_32_Re = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  out_results_32_Im = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  out_results_33_Re = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  out_results_33_Im = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  out_results_34_Re = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  out_results_34_Im = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  out_results_35_Re = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  out_results_35_Im = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  out_results_36_Re = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  out_results_36_Im = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  out_results_37_Re = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  out_results_37_Im = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  out_results_38_Re = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  out_results_38_Im = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  out_results_39_Re = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  out_results_39_Im = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  out_results_40_Re = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  out_results_40_Im = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  out_results_41_Re = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  out_results_41_Im = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  out_results_42_Re = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  out_results_42_Im = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  out_results_43_Re = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  out_results_43_Im = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  out_results_44_Re = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  out_results_44_Im = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  out_results_45_Re = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  out_results_45_Im = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  out_results_46_Re = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  out_results_46_Im = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  out_results_47_Re = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  out_results_47_Im = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  out_results_48_Re = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  out_results_48_Im = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  out_results_49_Re = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  out_results_49_Im = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  out_results_50_Re = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  out_results_50_Im = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  out_results_51_Re = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  out_results_51_Im = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  out_results_52_Re = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  out_results_52_Im = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  out_results_53_Re = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  out_results_53_Im = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  out_results_54_Re = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  out_results_54_Im = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  out_results_55_Re = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  out_results_55_Im = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  out_results_56_Re = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  out_results_56_Im = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  out_results_57_Re = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  out_results_57_Im = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  out_results_58_Re = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  out_results_58_Im = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  out_results_59_Re = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  out_results_59_Im = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  out_results_60_Re = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  out_results_60_Im = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  out_results_61_Re = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  out_results_61_Im = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  out_results_62_Re = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  out_results_62_Im = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  out_results_63_Re = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  out_results_63_Im = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  out_results_64_Re = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  out_results_64_Im = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  out_results_65_Re = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  out_results_65_Im = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  out_results_66_Re = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  out_results_66_Im = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  out_results_67_Re = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  out_results_67_Im = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  out_results_68_Re = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  out_results_68_Im = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  out_results_69_Re = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  out_results_69_Im = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  out_results_70_Re = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  out_results_70_Im = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  out_results_71_Re = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  out_results_71_Im = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  out_results_72_Re = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  out_results_72_Im = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  out_results_73_Re = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  out_results_73_Im = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  out_results_74_Re = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  out_results_74_Im = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  out_results_75_Re = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  out_results_75_Im = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  out_results_76_Re = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  out_results_76_Im = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  out_results_77_Re = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  out_results_77_Im = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  out_results_78_Re = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  out_results_78_Im = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  out_results_79_Re = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  out_results_79_Im = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  out_results_80_Re = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  out_results_80_Im = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  out_results_81_Re = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  out_results_81_Im = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  out_results_82_Re = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  out_results_82_Im = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  out_results_83_Re = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  out_results_83_Im = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  out_results_84_Re = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  out_results_84_Im = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  out_results_85_Re = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  out_results_85_Im = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  out_results_86_Re = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  out_results_86_Im = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  out_results_87_Re = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  out_results_87_Im = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  out_results_88_Re = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  out_results_88_Im = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  out_results_89_Re = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  out_results_89_Im = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  out_results_90_Re = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  out_results_90_Im = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  out_results_91_Re = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  out_results_91_Im = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  out_results_92_Re = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  out_results_92_Im = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  out_results_93_Re = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  out_results_93_Im = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  out_results_94_Re = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  out_results_94_Im = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  out_results_95_Re = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  out_results_95_Im = _RAND_209[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

