module cmplx_adj(
  input  [31:0] io_in_Re,
  input  [31:0] io_in_Im,
  input  [7:0]  io_in_adj,
  input         io_is_neg,
  input         io_is_flip,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  wire  sign_0 = io_in_Re[31]; // @[FFTDesigns.scala 4716:24]
  wire  sign_1 = io_in_Im[31]; // @[FFTDesigns.scala 4717:24]
  wire [7:0] exp_0 = io_in_Re[30:23]; // @[FFTDesigns.scala 4719:23]
  wire [7:0] exp_1 = io_in_Im[30:23]; // @[FFTDesigns.scala 4720:23]
  wire [22:0] frac_0 = io_in_Re[22:0]; // @[FFTDesigns.scala 4722:24]
  wire [22:0] frac_1 = io_in_Im[22:0]; // @[FFTDesigns.scala 4723:24]
  wire  new_sign_0 = io_is_neg ? ~sign_0 : sign_0; // @[FFTDesigns.scala 4725:20 4726:19 4729:19]
  wire  new_sign_1 = io_is_neg ? ~sign_1 : sign_1; // @[FFTDesigns.scala 4725:20 4727:19 4730:19]
  wire [7:0] _new_exp_0_T_1 = exp_0 - io_in_adj; // @[FFTDesigns.scala 4734:28]
  wire [7:0] new_exp_0 = exp_0 != 8'h0 ? _new_exp_0_T_1 : exp_0; // @[FFTDesigns.scala 4733:25 4734:18 4736:18]
  wire [7:0] _new_exp_1_T_1 = exp_1 - io_in_adj; // @[FFTDesigns.scala 4739:28]
  wire [7:0] new_exp_1 = exp_1 != 8'h0 ? _new_exp_1_T_1 : exp_1; // @[FFTDesigns.scala 4738:26 4739:18 4741:18]
  wire  _io_out_Re_T = ~new_sign_1; // @[FFTDesigns.scala 4745:21]
  wire [31:0] _io_out_Re_T_2 = {_io_out_Re_T,new_exp_1,frac_1}; // @[FFTDesigns.scala 4745:49]
  wire [31:0] _io_out_Im_T_1 = {new_sign_0,new_exp_0,frac_0}; // @[FFTDesigns.scala 4746:48]
  wire [31:0] _io_out_Im_T_3 = {new_sign_1,new_exp_1,frac_1}; // @[FFTDesigns.scala 4749:48]
  assign io_out_Re = io_is_flip ? _io_out_Re_T_2 : _io_out_Im_T_1; // @[FFTDesigns.scala 4744:21 4745:17 4748:17]
  assign io_out_Im = io_is_flip ? _io_out_Im_T_1 : _io_out_Im_T_3; // @[FFTDesigns.scala 4744:21 4746:17 4749:17]
endmodule
module full_subber(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[Arithmetic.scala 72:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[Arithmetic.scala 72:34]
  wire [8:0] result = _result_T_2[8:0]; // @[Arithmetic.scala 71:22 72:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 73:23]
  assign io_out_c = result[8]; // @[Arithmetic.scala 74:23]
endmodule
module twoscomplement(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _x_T = ~io_in; // @[Arithmetic.scala 28:16]
  assign io_out = 8'h1 + _x_T; // @[Arithmetic.scala 28:14]
endmodule
module full_adder(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 58:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 58:34]
  wire [24:0] result = _result_T_1[24:0]; // @[Arithmetic.scala 57:22 58:12]
  assign io_out_s = result[23:0]; // @[Arithmetic.scala 59:23]
  assign io_out_c = result[24]; // @[Arithmetic.scala 60:23]
endmodule
module twoscomplement_1(
  input  [23:0] io_in,
  output [23:0] io_out
);
  wire [23:0] _x_T = ~io_in; // @[Arithmetic.scala 28:16]
  assign io_out = 24'h1 + _x_T; // @[Arithmetic.scala 28:14]
endmodule
module shifter(
  input  [23:0] io_in_a,
  input  [4:0]  io_in_b,
  output [23:0] io_out_s
);
  wire [23:0] _result_T = io_in_a >> io_in_b; // @[Arithmetic.scala 42:25]
  wire [54:0] _GEN_0 = {{31'd0}, _result_T}; // @[Arithmetic.scala 41:26 42:14 44:14]
  assign io_out_s = _GEN_0[23:0]; // @[Arithmetic.scala 39:22]
endmodule
module leadingOneDetector(
  input  [23:0] io_in,
  output [4:0]  io_out
);
  wire [1:0] _hotValue_T = io_in[1] ? 2'h2 : 2'h1; // @[Mux.scala 47:70]
  wire [1:0] _hotValue_T_1 = io_in[2] ? 2'h3 : _hotValue_T; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_2 = io_in[3] ? 3'h4 : {{1'd0}, _hotValue_T_1}; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_3 = io_in[4] ? 3'h5 : _hotValue_T_2; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_4 = io_in[5] ? 3'h6 : _hotValue_T_3; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_5 = io_in[6] ? 3'h7 : _hotValue_T_4; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_6 = io_in[7] ? 4'h8 : {{1'd0}, _hotValue_T_5}; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_7 = io_in[8] ? 4'h9 : _hotValue_T_6; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_8 = io_in[9] ? 4'ha : _hotValue_T_7; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_9 = io_in[10] ? 4'hb : _hotValue_T_8; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_10 = io_in[11] ? 4'hc : _hotValue_T_9; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_11 = io_in[12] ? 4'hd : _hotValue_T_10; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_12 = io_in[13] ? 4'he : _hotValue_T_11; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_13 = io_in[14] ? 4'hf : _hotValue_T_12; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_14 = io_in[15] ? 5'h10 : {{1'd0}, _hotValue_T_13}; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_15 = io_in[16] ? 5'h11 : _hotValue_T_14; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_16 = io_in[17] ? 5'h12 : _hotValue_T_15; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_17 = io_in[18] ? 5'h13 : _hotValue_T_16; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_18 = io_in[19] ? 5'h14 : _hotValue_T_17; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_19 = io_in[20] ? 5'h15 : _hotValue_T_18; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_20 = io_in[21] ? 5'h16 : _hotValue_T_19; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_21 = io_in[22] ? 5'h17 : _hotValue_T_20; // @[Mux.scala 47:70]
  assign io_out = io_in[23] ? 5'h18 : _hotValue_T_21; // @[Mux.scala 47:70]
endmodule
module FP_adder(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 76:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 76:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 76:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 76:24]
  wire [7:0] complement_io_in; // @[FPArithmetic.scala 82:28]
  wire [7:0] complement_io_out; // @[FPArithmetic.scala 82:28]
  wire [23:0] adder_io_in_a; // @[FPArithmetic.scala 86:23]
  wire [23:0] adder_io_in_b; // @[FPArithmetic.scala 86:23]
  wire [23:0] adder_io_out_s; // @[FPArithmetic.scala 86:23]
  wire  adder_io_out_c; // @[FPArithmetic.scala 86:23]
  wire [23:0] complementN_0_io_in; // @[FPArithmetic.scala 92:31]
  wire [23:0] complementN_0_io_out; // @[FPArithmetic.scala 92:31]
  wire [23:0] complementN_1_io_in; // @[FPArithmetic.scala 94:31]
  wire [23:0] complementN_1_io_out; // @[FPArithmetic.scala 94:31]
  wire [23:0] shifter_io_in_a; // @[FPArithmetic.scala 98:25]
  wire [4:0] shifter_io_in_b; // @[FPArithmetic.scala 98:25]
  wire [23:0] shifter_io_out_s; // @[FPArithmetic.scala 98:25]
  wire [23:0] complementN_2_io_in; // @[FPArithmetic.scala 143:31]
  wire [23:0] complementN_2_io_out; // @[FPArithmetic.scala 143:31]
  wire [23:0] leadingOneFinder_io_in; // @[FPArithmetic.scala 163:34]
  wire [4:0] leadingOneFinder_io_out; // @[FPArithmetic.scala 163:34]
  wire [7:0] subber2_io_in_a; // @[FPArithmetic.scala 165:25]
  wire [7:0] subber2_io_in_b; // @[FPArithmetic.scala 165:25]
  wire [7:0] subber2_io_out_s; // @[FPArithmetic.scala 165:25]
  wire  subber2_io_out_c; // @[FPArithmetic.scala 165:25]
  wire  sign_0 = io_in_a[31]; // @[FPArithmetic.scala 38:23]
  wire  sign_1 = io_in_b[31]; // @[FPArithmetic.scala 39:23]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 43:62]
  wire [8:0] _GEN_31 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 43:34]
  wire [8:0] _GEN_0 = _GEN_31 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 43:68 44:14 46:14]
  wire [8:0] _GEN_32 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 48:34]
  wire [8:0] _GEN_1 = _GEN_32 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 48:68 49:14 51:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 56:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 57:23]
  wire [23:0] whole_frac_0 = {1'h1,frac_0}; // @[FPArithmetic.scala 61:26]
  wire [23:0] whole_frac_1 = {1'h1,frac_1}; // @[FPArithmetic.scala 62:26]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 42:19]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 42:19]
  wire [7:0] out_exp = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 104:34 105:15 115:15]
  wire [7:0] sub_exp = subber_io_out_c ? complement_io_out : subber_io_out_s; // @[FPArithmetic.scala 104:34 106:15 116:15]
  wire  out_s = subber_io_out_c ? sign_1 : sign_0; // @[FPArithmetic.scala 104:34 107:13 117:13]
  wire [22:0] out_frac = subber_io_out_c ? frac_1 : frac_0; // @[FPArithmetic.scala 104:34 108:16 118:16]
  wire [23:0] _GEN_8 = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 104:34 112:21 87:19]
  wire [23:0] _GEN_9 = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 104:34 88:19 122:21]
  wire  _new_s_T = ~adder_io_out_c; // @[FPArithmetic.scala 138:15]
  wire  _D_T_1 = sign_0 ^ sign_1; // @[FPArithmetic.scala 151:39]
  wire  D = _new_s_T | sign_0 ^ sign_1; // @[FPArithmetic.scala 151:28]
  wire  E = _new_s_T & ~adder_io_out_s[23] | _new_s_T & ~_D_T_1 | adder_io_out_c & adder_io_out_s[23] & _D_T_1; // @[FPArithmetic.scala 154:99]
  wire  _GEN_25 = sub_exp >= 8'h17 ? out_s : ~adder_io_out_c & sign_0 | sign_0 & sign_1 | ~adder_io_out_c & sign_1; // @[FPArithmetic.scala 138:11 173:39 174:13]
  wire  new_s = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 1'h0 : _GEN_25; // @[FPArithmetic.scala 169:62 170:13]
  wire [23:0] adder_result = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 157:18 158:47 159:20]
  wire [4:0] _subber2_io_in_b_T_1 = 5'h18 - leadingOneFinder_io_out; // @[FPArithmetic.scala 167:42]
  wire [8:0] _GEN_33 = {{1'd0}, out_exp}; // @[FPArithmetic.scala 181:20]
  wire [23:0] _new_out_frac_T_2 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 183:51]
  wire [7:0] _new_out_exp_T_3 = out_exp + 8'h1; // @[FPArithmetic.scala 185:32]
  wire [8:0] _GEN_13 = _GEN_33 == _T_2 ? _T_2 : {{1'd0}, _new_out_exp_T_3}; // @[FPArithmetic.scala 181:56 182:21 185:21]
  wire [23:0] _GEN_14 = _GEN_33 == _T_2 ? _new_out_frac_T_2 : {{1'd0}, adder_result[23:1]}; // @[FPArithmetic.scala 181:56 183:22 186:22]
  wire [53:0] _GEN_2 = {{31'd0}, adder_result[22:0]}; // @[FPArithmetic.scala 197:57]
  wire [53:0] _new_out_frac_T_7 = _GEN_2 << _subber2_io_in_b_T_1; // @[FPArithmetic.scala 197:57]
  wire [7:0] _GEN_15 = subber2_io_out_c ? 8'h1 : subber2_io_out_s; // @[FPArithmetic.scala 192:39 193:23 196:23]
  wire [53:0] _GEN_16 = subber2_io_out_c ? 54'h400000 : _new_out_frac_T_7; // @[FPArithmetic.scala 192:39 194:24 197:24]
  wire [7:0] _GEN_17 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:0
    ]) ? 8'h0 : _GEN_15; // @[FPArithmetic.scala 189:141 190:21]
  wire [53:0] _GEN_18 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:
    0]) ? 54'h0 : _GEN_16; // @[FPArithmetic.scala 189:141 139:18]
  wire [7:0] _GEN_19 = D ? _GEN_17 : 8'h0; // @[FPArithmetic.scala 140:17 188:26]
  wire [53:0] _GEN_20 = D ? _GEN_18 : 54'h0; // @[FPArithmetic.scala 139:18 188:26]
  wire [8:0] _GEN_21 = ~D ? _GEN_13 : {{1'd0}, _GEN_19}; // @[FPArithmetic.scala 180:26]
  wire [53:0] _GEN_22 = ~D ? {{30'd0}, _GEN_14} : _GEN_20; // @[FPArithmetic.scala 180:26]
  wire [8:0] _GEN_23 = E ? {{1'd0}, out_exp} : _GEN_21; // @[FPArithmetic.scala 177:26 178:19]
  wire [53:0] _GEN_24 = E ? {{31'd0}, adder_result[22:0]} : _GEN_22; // @[FPArithmetic.scala 177:26 179:20]
  wire [53:0] _GEN_26 = sub_exp >= 8'h17 ? {{31'd0}, out_frac} : _GEN_24; // @[FPArithmetic.scala 173:39 175:20]
  wire [8:0] _GEN_27 = sub_exp >= 8'h17 ? {{1'd0}, out_exp} : _GEN_23; // @[FPArithmetic.scala 173:39 176:19]
  wire [8:0] _GEN_29 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 9'h0 : _GEN_27; // @[FPArithmetic.scala 169:62 171:19]
  wire [53:0] _GEN_30 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 54'h0 : _GEN_26; // @[FPArithmetic.scala 169:62 172:20]
  reg [31:0] reg_out_s; // @[FPArithmetic.scala 201:28]
  wire [7:0] new_out_exp = _GEN_29[7:0]; // @[FPArithmetic.scala 137:27]
  wire [22:0] new_out_frac = _GEN_30[22:0]; // @[FPArithmetic.scala 136:28]
  wire [31:0] _reg_out_s_T_1 = {new_s,new_out_exp,new_out_frac}; // @[FPArithmetic.scala 203:39]
  full_subber subber ( // @[FPArithmetic.scala 76:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complement ( // @[FPArithmetic.scala 82:28]
    .io_in(complement_io_in),
    .io_out(complement_io_out)
  );
  full_adder adder ( // @[FPArithmetic.scala 86:23]
    .io_in_a(adder_io_in_a),
    .io_in_b(adder_io_in_b),
    .io_out_s(adder_io_out_s),
    .io_out_c(adder_io_out_c)
  );
  twoscomplement_1 complementN_0 ( // @[FPArithmetic.scala 92:31]
    .io_in(complementN_0_io_in),
    .io_out(complementN_0_io_out)
  );
  twoscomplement_1 complementN_1 ( // @[FPArithmetic.scala 94:31]
    .io_in(complementN_1_io_in),
    .io_out(complementN_1_io_out)
  );
  shifter shifter ( // @[FPArithmetic.scala 98:25]
    .io_in_a(shifter_io_in_a),
    .io_in_b(shifter_io_in_b),
    .io_out_s(shifter_io_out_s)
  );
  twoscomplement_1 complementN_2 ( // @[FPArithmetic.scala 143:31]
    .io_in(complementN_2_io_in),
    .io_out(complementN_2_io_out)
  );
  leadingOneDetector leadingOneFinder ( // @[FPArithmetic.scala 163:34]
    .io_in(leadingOneFinder_io_in),
    .io_out(leadingOneFinder_io_out)
  );
  full_subber subber2 ( // @[FPArithmetic.scala 165:25]
    .io_in_a(subber2_io_in_a),
    .io_in_b(subber2_io_in_b),
    .io_out_s(subber2_io_out_s),
    .io_out_c(subber2_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FPArithmetic.scala 205:14]
  assign subber_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 42:19]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 42:19]
  assign complement_io_in = subber_io_out_s; // @[FPArithmetic.scala 83:22]
  assign adder_io_in_a = sign_0 & ~sign_1 ? complementN_0_io_out : _GEN_8; // @[FPArithmetic.scala 127:45 128:21]
  assign adder_io_in_b = sign_1 & ~sign_0 ? complementN_1_io_out : _GEN_9; // @[FPArithmetic.scala 131:45 132:21]
  assign complementN_0_io_in = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 104:34 112:21 87:19]
  assign complementN_1_io_in = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 104:34 88:19 122:21]
  assign shifter_io_in_a = subber_io_out_c ? whole_frac_0 : whole_frac_1; // @[FPArithmetic.scala 104:34 109:23 119:23]
  assign shifter_io_in_b = sub_exp[4:0];
  assign complementN_2_io_in = adder_io_out_s; // @[FPArithmetic.scala 144:25]
  assign leadingOneFinder_io_in = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 157:18 158:47 159:20]
  assign subber2_io_in_a = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 104:34 105:15 115:15]
  assign subber2_io_in_b = {{3'd0}, _subber2_io_in_b_T_1}; // @[FPArithmetic.scala 167:21]
  always @(posedge clock) begin
    if (reset) begin // @[FPArithmetic.scala 201:28]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 201:28]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FPArithmetic.scala 203:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_out_s = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexAdder(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_adder_clock; // @[FPComplex.scala 21:25]
  wire  FP_adder_reset; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 21:25]
  wire  FP_adder_1_clock; // @[FPComplex.scala 21:25]
  wire  FP_adder_1_reset; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_in_a; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_in_b; // @[FPComplex.scala 21:25]
  wire [31:0] FP_adder_1_io_out_s; // @[FPComplex.scala 21:25]
  FP_adder FP_adder ( // @[FPComplex.scala 21:25]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_adder FP_adder_1 ( // @[FPComplex.scala 21:25]
    .clock(FP_adder_1_clock),
    .reset(FP_adder_1_reset),
    .io_in_a(FP_adder_1_io_in_a),
    .io_in_b(FP_adder_1_io_in_b),
    .io_out_s(FP_adder_1_io_out_s)
  );
  assign io_out_s_Re = FP_adder_io_out_s; // @[FPComplex.scala 28:17]
  assign io_out_s_Im = FP_adder_1_io_out_s; // @[FPComplex.scala 29:17]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = io_in_a_Re; // @[FPComplex.scala 24:23]
  assign FP_adder_io_in_b = io_in_b_Re; // @[FPComplex.scala 25:23]
  assign FP_adder_1_clock = clock;
  assign FP_adder_1_reset = reset;
  assign FP_adder_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 26:23]
  assign FP_adder_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 27:23]
endmodule
module FPComplexMultiAdder(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  wire  FPComplexAdder_clock; // @[FPComplex.scala 524:30]
  wire  FPComplexAdder_reset; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_in_a_Re; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_in_a_Im; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_in_b_Re; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_in_b_Im; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_out_s_Re; // @[FPComplex.scala 524:30]
  wire [31:0] FPComplexAdder_io_out_s_Im; // @[FPComplex.scala 524:30]
  FPComplexAdder FPComplexAdder ( // @[FPComplex.scala 524:30]
    .clock(FPComplexAdder_clock),
    .reset(FPComplexAdder_reset),
    .io_in_a_Re(FPComplexAdder_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_io_out_s_Im)
  );
  assign io_out_Re = FPComplexAdder_io_out_s_Re; // @[FPComplex.scala 642:16]
  assign io_out_Im = FPComplexAdder_io_out_s_Im; // @[FPComplex.scala 642:16]
  assign FPComplexAdder_clock = clock;
  assign FPComplexAdder_reset = reset;
  assign FPComplexAdder_io_in_a_Re = io_in_0_Re; // @[FPComplex.scala 604:42]
  assign FPComplexAdder_io_in_a_Im = io_in_0_Im; // @[FPComplex.scala 604:42]
  assign FPComplexAdder_io_in_b_Re = io_in_1_Re; // @[FPComplex.scala 605:42]
  assign FPComplexAdder_io_in_b_Im = io_in_1_Im; // @[FPComplex.scala 605:42]
endmodule
module DFT_r_V1_nonregout(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im
);
  wire [31:0] cmplx_adj_io_in_Re; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_in_Im; // @[FFTDesigns.scala 1808:22]
  wire [7:0] cmplx_adj_io_in_adj; // @[FFTDesigns.scala 1808:22]
  wire  cmplx_adj_io_is_neg; // @[FFTDesigns.scala 1808:22]
  wire  cmplx_adj_io_is_flip; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_out_Re; // @[FFTDesigns.scala 1808:22]
  wire [31:0] cmplx_adj_io_out_Im; // @[FFTDesigns.scala 1808:22]
  wire  FPComplexMultiAdder_clock; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_reset; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_0_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_0_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_1_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_in_1_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_1_clock; // @[FFTDesigns.scala 1839:26]
  wire  FPComplexMultiAdder_1_reset; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_1_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_in_1_Im; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 1839:26]
  wire [31:0] FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 1839:26]
  cmplx_adj cmplx_adj ( // @[FFTDesigns.scala 1808:22]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder ( // @[FFTDesigns.scala 1839:26]
    .clock(FPComplexMultiAdder_clock),
    .reset(FPComplexMultiAdder_reset),
    .io_in_0_Re(FPComplexMultiAdder_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_io_in_1_Im),
    .io_out_Re(FPComplexMultiAdder_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_io_out_Im)
  );
  FPComplexMultiAdder FPComplexMultiAdder_1 ( // @[FFTDesigns.scala 1839:26]
    .clock(FPComplexMultiAdder_1_clock),
    .reset(FPComplexMultiAdder_1_reset),
    .io_in_0_Re(FPComplexMultiAdder_1_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_1_io_in_0_Im),
    .io_in_1_Re(FPComplexMultiAdder_1_io_in_1_Re),
    .io_in_1_Im(FPComplexMultiAdder_1_io_in_1_Im),
    .io_out_Re(FPComplexMultiAdder_1_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_1_io_out_Im)
  );
  assign io_out_0_Re = FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 1911:17]
  assign io_out_0_Im = FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 1911:17]
  assign io_out_1_Re = FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 1911:17]
  assign io_out_1_Im = FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 1911:17]
  assign cmplx_adj_io_in_Re = io_in_1_Re; // @[FFTDesigns.scala 1820:27]
  assign cmplx_adj_io_in_Im = io_in_1_Im; // @[FFTDesigns.scala 1820:27]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FFTDesigns.scala 1821:31]
  assign cmplx_adj_io_is_neg = 1'h1; // @[FFTDesigns.scala 1822:31]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FFTDesigns.scala 1823:32]
  assign FPComplexMultiAdder_clock = clock;
  assign FPComplexMultiAdder_reset = reset;
  assign FPComplexMultiAdder_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 1891:30]
  assign FPComplexMultiAdder_1_clock = clock;
  assign FPComplexMultiAdder_1_reset = reset;
  assign FPComplexMultiAdder_1_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 1896:32]
  assign FPComplexMultiAdder_1_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 1896:32]
  assign FPComplexMultiAdder_1_io_in_1_Re = cmplx_adj_io_out_Re; // @[FFTDesigns.scala 1818:24 1824:42]
  assign FPComplexMultiAdder_1_io_in_1_Im = cmplx_adj_io_out_Im; // @[FFTDesigns.scala 1818:24 1824:42]
endmodule
module DFT_r_v2(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im
);
  wire  DFT_r_V1_nonregout_clock; // @[FFTDesigns.scala 169:24]
  wire  DFT_r_V1_nonregout_reset; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_0_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_0_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_1_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_in_1_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_0_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_0_Im; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_1_Re; // @[FFTDesigns.scala 169:24]
  wire [31:0] DFT_r_V1_nonregout_io_out_1_Im; // @[FFTDesigns.scala 169:24]
  DFT_r_V1_nonregout DFT_r_V1_nonregout ( // @[FFTDesigns.scala 169:24]
    .clock(DFT_r_V1_nonregout_clock),
    .reset(DFT_r_V1_nonregout_reset),
    .io_in_0_Re(DFT_r_V1_nonregout_io_in_0_Re),
    .io_in_0_Im(DFT_r_V1_nonregout_io_in_0_Im),
    .io_in_1_Re(DFT_r_V1_nonregout_io_in_1_Re),
    .io_in_1_Im(DFT_r_V1_nonregout_io_in_1_Im),
    .io_out_0_Re(DFT_r_V1_nonregout_io_out_0_Re),
    .io_out_0_Im(DFT_r_V1_nonregout_io_out_0_Im),
    .io_out_1_Re(DFT_r_V1_nonregout_io_out_1_Re),
    .io_out_1_Im(DFT_r_V1_nonregout_io_out_1_Im)
  );
  assign io_out_0_Re = DFT_r_V1_nonregout_io_out_0_Re; // @[FFTDesigns.scala 171:14]
  assign io_out_0_Im = DFT_r_V1_nonregout_io_out_0_Im; // @[FFTDesigns.scala 171:14]
  assign io_out_1_Re = DFT_r_V1_nonregout_io_out_1_Re; // @[FFTDesigns.scala 171:14]
  assign io_out_1_Im = DFT_r_V1_nonregout_io_out_1_Im; // @[FFTDesigns.scala 171:14]
  assign DFT_r_V1_nonregout_clock = clock;
  assign DFT_r_V1_nonregout_reset = reset;
  assign DFT_r_V1_nonregout_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 170:15]
  assign DFT_r_V1_nonregout_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 170:15]
endmodule
module RAM_Block(
  input         clock,
  input  [1:0]  io_in_raddr,
  input  [1:0]  io_in_waddr,
  input  [31:0] io_in_data_Re,
  input  [31:0] io_in_data_Im,
  input         io_re,
  input         io_wr,
  input         io_en,
  output [31:0] io_out_data_Re,
  output [31:0] io_out_data_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_0_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Im; // @[FFTDesigns.scala 3286:18]
  wire [31:0] _GEN_17 = 2'h1 == io_in_raddr ? mem_1_Im : mem_0_Im; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_18 = 2'h2 == io_in_raddr ? mem_2_Im : _GEN_17; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_19 = 2'h3 == io_in_raddr ? mem_3_Im : _GEN_18; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_21 = 2'h1 == io_in_raddr ? mem_1_Re : mem_0_Re; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_22 = 2'h2 == io_in_raddr ? mem_2_Re : _GEN_21; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_23 = 2'h3 == io_in_raddr ? mem_3_Re : _GEN_22; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_24 = io_re ? _GEN_19 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3295:24]
  wire [31:0] _GEN_25 = io_re ? _GEN_23 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3294:24]
  assign io_out_data_Re = io_en ? _GEN_25 : 32'h0; // @[FFTDesigns.scala 3287:16 3298:22]
  assign io_out_data_Im = io_en ? _GEN_24 : 32'h0; // @[FFTDesigns.scala 3287:16 3299:22]
  always @(posedge clock) begin
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (2'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (2'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (2'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (2'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (2'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (2'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (2'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (2'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_3_Im = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PermutationModuleStreamed(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [3:0]  io_in_config_0,
  input  [3:0]  io_in_config_1,
  input  [3:0]  io_in_config_2,
  input  [3:0]  io_in_config_3,
  input  [3:0]  io_in_config_4,
  input  [3:0]  io_in_config_5,
  input  [3:0]  io_in_config_6,
  input  [3:0]  io_in_config_7,
  input  [3:0]  io_in_config_8,
  input  [3:0]  io_in_config_9,
  input  [3:0]  io_in_config_10,
  input  [3:0]  io_in_config_11,
  input  [3:0]  io_in_config_12,
  input  [3:0]  io_in_config_13,
  input  [3:0]  io_in_config_14,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
  wire  _T = io_in_config_0 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_1 = io_in_config_1 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_2 = io_in_config_2 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_3 = io_in_config_3 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_4 = io_in_config_4 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_5 = io_in_config_5 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_6 = io_in_config_6 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_7 = io_in_config_7 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_8 = io_in_config_8 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_9 = io_in_config_9 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_10 = io_in_config_10 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_11 = io_in_config_11 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_12 = io_in_config_12 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_13 = io_in_config_13 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_14 = io_in_config_14 == 4'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_16 = io_in_config_0 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_17 = io_in_config_1 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_18 = io_in_config_2 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_19 = io_in_config_3 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_20 = io_in_config_4 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_21 = io_in_config_5 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_22 = io_in_config_6 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_23 = io_in_config_7 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_24 = io_in_config_8 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_25 = io_in_config_9 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_26 = io_in_config_10 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_27 = io_in_config_11 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_28 = io_in_config_12 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_29 = io_in_config_13 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_30 = io_in_config_14 == 4'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_32 = io_in_config_0 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_33 = io_in_config_1 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_34 = io_in_config_2 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_35 = io_in_config_3 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_36 = io_in_config_4 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_37 = io_in_config_5 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_38 = io_in_config_6 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_39 = io_in_config_7 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_40 = io_in_config_8 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_41 = io_in_config_9 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_42 = io_in_config_10 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_43 = io_in_config_11 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_44 = io_in_config_12 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_45 = io_in_config_13 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_46 = io_in_config_14 == 4'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_48 = io_in_config_0 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_49 = io_in_config_1 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_50 = io_in_config_2 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_51 = io_in_config_3 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_52 = io_in_config_4 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_53 = io_in_config_5 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_54 = io_in_config_6 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_55 = io_in_config_7 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_56 = io_in_config_8 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_57 = io_in_config_9 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_58 = io_in_config_10 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_59 = io_in_config_11 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_60 = io_in_config_12 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_61 = io_in_config_13 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_62 = io_in_config_14 == 4'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_64 = io_in_config_0 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_65 = io_in_config_1 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_66 = io_in_config_2 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_67 = io_in_config_3 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_68 = io_in_config_4 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_69 = io_in_config_5 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_70 = io_in_config_6 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_71 = io_in_config_7 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_72 = io_in_config_8 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_73 = io_in_config_9 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_74 = io_in_config_10 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_75 = io_in_config_11 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_76 = io_in_config_12 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_77 = io_in_config_13 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_78 = io_in_config_14 == 4'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_80 = io_in_config_0 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_81 = io_in_config_1 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_82 = io_in_config_2 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_83 = io_in_config_3 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_84 = io_in_config_4 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_85 = io_in_config_5 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_86 = io_in_config_6 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_87 = io_in_config_7 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_88 = io_in_config_8 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_89 = io_in_config_9 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_90 = io_in_config_10 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_91 = io_in_config_11 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_92 = io_in_config_12 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_93 = io_in_config_13 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_94 = io_in_config_14 == 4'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_96 = io_in_config_0 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_97 = io_in_config_1 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_98 = io_in_config_2 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_99 = io_in_config_3 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_100 = io_in_config_4 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_101 = io_in_config_5 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_102 = io_in_config_6 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_103 = io_in_config_7 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_104 = io_in_config_8 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_105 = io_in_config_9 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_106 = io_in_config_10 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_107 = io_in_config_11 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_108 = io_in_config_12 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_109 = io_in_config_13 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_110 = io_in_config_14 == 4'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_112 = io_in_config_0 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_113 = io_in_config_1 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_114 = io_in_config_2 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_115 = io_in_config_3 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_116 = io_in_config_4 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_117 = io_in_config_5 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_118 = io_in_config_6 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_119 = io_in_config_7 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_120 = io_in_config_8 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_121 = io_in_config_9 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_122 = io_in_config_10 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_123 = io_in_config_11 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_124 = io_in_config_12 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_125 = io_in_config_13 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_126 = io_in_config_14 == 4'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_128 = io_in_config_0 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_129 = io_in_config_1 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_130 = io_in_config_2 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_131 = io_in_config_3 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_132 = io_in_config_4 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_133 = io_in_config_5 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_134 = io_in_config_6 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_135 = io_in_config_7 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_136 = io_in_config_8 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_137 = io_in_config_9 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_138 = io_in_config_10 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_139 = io_in_config_11 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_140 = io_in_config_12 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_141 = io_in_config_13 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_142 = io_in_config_14 == 4'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_144 = io_in_config_0 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_145 = io_in_config_1 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_146 = io_in_config_2 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_147 = io_in_config_3 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_148 = io_in_config_4 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_149 = io_in_config_5 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_150 = io_in_config_6 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_151 = io_in_config_7 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_152 = io_in_config_8 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_153 = io_in_config_9 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_154 = io_in_config_10 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_155 = io_in_config_11 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_156 = io_in_config_12 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_157 = io_in_config_13 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_158 = io_in_config_14 == 4'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_160 = io_in_config_0 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_161 = io_in_config_1 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_162 = io_in_config_2 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_163 = io_in_config_3 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_164 = io_in_config_4 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_165 = io_in_config_5 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_166 = io_in_config_6 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_167 = io_in_config_7 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_168 = io_in_config_8 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_169 = io_in_config_9 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_170 = io_in_config_10 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_171 = io_in_config_11 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_172 = io_in_config_12 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_173 = io_in_config_13 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_174 = io_in_config_14 == 4'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_176 = io_in_config_0 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_177 = io_in_config_1 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_178 = io_in_config_2 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_179 = io_in_config_3 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_180 = io_in_config_4 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_181 = io_in_config_5 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_182 = io_in_config_6 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_183 = io_in_config_7 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_184 = io_in_config_8 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_185 = io_in_config_9 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_186 = io_in_config_10 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_187 = io_in_config_11 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_188 = io_in_config_12 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_189 = io_in_config_13 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_190 = io_in_config_14 == 4'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_192 = io_in_config_0 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_193 = io_in_config_1 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_194 = io_in_config_2 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_195 = io_in_config_3 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_196 = io_in_config_4 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_197 = io_in_config_5 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_198 = io_in_config_6 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_199 = io_in_config_7 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_200 = io_in_config_8 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_201 = io_in_config_9 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_202 = io_in_config_10 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_203 = io_in_config_11 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_204 = io_in_config_12 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_205 = io_in_config_13 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_206 = io_in_config_14 == 4'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_208 = io_in_config_0 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_209 = io_in_config_1 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_210 = io_in_config_2 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_211 = io_in_config_3 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_212 = io_in_config_4 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_213 = io_in_config_5 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_214 = io_in_config_6 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_215 = io_in_config_7 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_216 = io_in_config_8 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_217 = io_in_config_9 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_218 = io_in_config_10 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_219 = io_in_config_11 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_220 = io_in_config_12 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_221 = io_in_config_13 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_222 = io_in_config_14 == 4'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_224 = io_in_config_0 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_225 = io_in_config_1 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_226 = io_in_config_2 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_227 = io_in_config_3 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_228 = io_in_config_4 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_229 = io_in_config_5 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_230 = io_in_config_6 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_231 = io_in_config_7 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_232 = io_in_config_8 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_233 = io_in_config_9 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_234 = io_in_config_10 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_235 = io_in_config_11 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_236 = io_in_config_12 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_237 = io_in_config_13 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_238 = io_in_config_14 == 4'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_240 = io_in_config_0 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_241 = io_in_config_1 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_242 = io_in_config_2 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_243 = io_in_config_3 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_244 = io_in_config_4 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_245 = io_in_config_5 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_246 = io_in_config_6 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_247 = io_in_config_7 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_248 = io_in_config_8 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_249 = io_in_config_9 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_250 = io_in_config_10 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_251 = io_in_config_11 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_252 = io_in_config_12 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_253 = io_in_config_13 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_254 = io_in_config_14 == 4'hf; // @[FFTDesigns.scala 3194:35]
  wire [3:0] _pms_pmx_T = _T_14 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_1 = _T_13 ? 4'hd : _pms_pmx_T; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_2 = _T_12 ? 4'hc : _pms_pmx_T_1; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_3 = _T_11 ? 4'hb : _pms_pmx_T_2; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_4 = _T_10 ? 4'ha : _pms_pmx_T_3; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_5 = _T_9 ? 4'h9 : _pms_pmx_T_4; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_6 = _T_8 ? 4'h8 : _pms_pmx_T_5; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_7 = _T_7 ? 4'h7 : _pms_pmx_T_6; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_8 = _T_6 ? 4'h6 : _pms_pmx_T_7; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_9 = _T_5 ? 4'h5 : _pms_pmx_T_8; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_10 = _T_4 ? 4'h4 : _pms_pmx_T_9; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_11 = _T_3 ? 4'h3 : _pms_pmx_T_10; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_12 = _T_2 ? 4'h2 : _pms_pmx_T_11; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_13 = _T_1 ? 4'h1 : _pms_pmx_T_12; // @[Mux.scala 47:70]
  wire [3:0] pms_0 = _T ? 4'h0 : _pms_pmx_T_13; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_14 = _T_30 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_15 = _T_29 ? 4'hd : _pms_pmx_T_14; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_16 = _T_28 ? 4'hc : _pms_pmx_T_15; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_17 = _T_27 ? 4'hb : _pms_pmx_T_16; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_18 = _T_26 ? 4'ha : _pms_pmx_T_17; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_19 = _T_25 ? 4'h9 : _pms_pmx_T_18; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_20 = _T_24 ? 4'h8 : _pms_pmx_T_19; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_21 = _T_23 ? 4'h7 : _pms_pmx_T_20; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_22 = _T_22 ? 4'h6 : _pms_pmx_T_21; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_23 = _T_21 ? 4'h5 : _pms_pmx_T_22; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_24 = _T_20 ? 4'h4 : _pms_pmx_T_23; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_25 = _T_19 ? 4'h3 : _pms_pmx_T_24; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_26 = _T_18 ? 4'h2 : _pms_pmx_T_25; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_27 = _T_17 ? 4'h1 : _pms_pmx_T_26; // @[Mux.scala 47:70]
  wire [3:0] pms_1 = _T_16 ? 4'h0 : _pms_pmx_T_27; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_28 = _T_46 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_29 = _T_45 ? 4'hd : _pms_pmx_T_28; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_30 = _T_44 ? 4'hc : _pms_pmx_T_29; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_31 = _T_43 ? 4'hb : _pms_pmx_T_30; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_32 = _T_42 ? 4'ha : _pms_pmx_T_31; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_33 = _T_41 ? 4'h9 : _pms_pmx_T_32; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_34 = _T_40 ? 4'h8 : _pms_pmx_T_33; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_35 = _T_39 ? 4'h7 : _pms_pmx_T_34; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_36 = _T_38 ? 4'h6 : _pms_pmx_T_35; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_37 = _T_37 ? 4'h5 : _pms_pmx_T_36; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_38 = _T_36 ? 4'h4 : _pms_pmx_T_37; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_39 = _T_35 ? 4'h3 : _pms_pmx_T_38; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_40 = _T_34 ? 4'h2 : _pms_pmx_T_39; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_41 = _T_33 ? 4'h1 : _pms_pmx_T_40; // @[Mux.scala 47:70]
  wire [3:0] pms_2 = _T_32 ? 4'h0 : _pms_pmx_T_41; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_42 = _T_62 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_43 = _T_61 ? 4'hd : _pms_pmx_T_42; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_44 = _T_60 ? 4'hc : _pms_pmx_T_43; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_45 = _T_59 ? 4'hb : _pms_pmx_T_44; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_46 = _T_58 ? 4'ha : _pms_pmx_T_45; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_47 = _T_57 ? 4'h9 : _pms_pmx_T_46; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_48 = _T_56 ? 4'h8 : _pms_pmx_T_47; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_49 = _T_55 ? 4'h7 : _pms_pmx_T_48; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_50 = _T_54 ? 4'h6 : _pms_pmx_T_49; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_51 = _T_53 ? 4'h5 : _pms_pmx_T_50; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_52 = _T_52 ? 4'h4 : _pms_pmx_T_51; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_53 = _T_51 ? 4'h3 : _pms_pmx_T_52; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_54 = _T_50 ? 4'h2 : _pms_pmx_T_53; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_55 = _T_49 ? 4'h1 : _pms_pmx_T_54; // @[Mux.scala 47:70]
  wire [3:0] pms_3 = _T_48 ? 4'h0 : _pms_pmx_T_55; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_56 = _T_78 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_57 = _T_77 ? 4'hd : _pms_pmx_T_56; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_58 = _T_76 ? 4'hc : _pms_pmx_T_57; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_59 = _T_75 ? 4'hb : _pms_pmx_T_58; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_60 = _T_74 ? 4'ha : _pms_pmx_T_59; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_61 = _T_73 ? 4'h9 : _pms_pmx_T_60; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_62 = _T_72 ? 4'h8 : _pms_pmx_T_61; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_63 = _T_71 ? 4'h7 : _pms_pmx_T_62; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_64 = _T_70 ? 4'h6 : _pms_pmx_T_63; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_65 = _T_69 ? 4'h5 : _pms_pmx_T_64; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_66 = _T_68 ? 4'h4 : _pms_pmx_T_65; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_67 = _T_67 ? 4'h3 : _pms_pmx_T_66; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_68 = _T_66 ? 4'h2 : _pms_pmx_T_67; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_69 = _T_65 ? 4'h1 : _pms_pmx_T_68; // @[Mux.scala 47:70]
  wire [3:0] pms_4 = _T_64 ? 4'h0 : _pms_pmx_T_69; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_70 = _T_94 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_71 = _T_93 ? 4'hd : _pms_pmx_T_70; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_72 = _T_92 ? 4'hc : _pms_pmx_T_71; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_73 = _T_91 ? 4'hb : _pms_pmx_T_72; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_74 = _T_90 ? 4'ha : _pms_pmx_T_73; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_75 = _T_89 ? 4'h9 : _pms_pmx_T_74; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_76 = _T_88 ? 4'h8 : _pms_pmx_T_75; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_77 = _T_87 ? 4'h7 : _pms_pmx_T_76; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_78 = _T_86 ? 4'h6 : _pms_pmx_T_77; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_79 = _T_85 ? 4'h5 : _pms_pmx_T_78; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_80 = _T_84 ? 4'h4 : _pms_pmx_T_79; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_81 = _T_83 ? 4'h3 : _pms_pmx_T_80; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_82 = _T_82 ? 4'h2 : _pms_pmx_T_81; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_83 = _T_81 ? 4'h1 : _pms_pmx_T_82; // @[Mux.scala 47:70]
  wire [3:0] pms_5 = _T_80 ? 4'h0 : _pms_pmx_T_83; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_84 = _T_110 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_85 = _T_109 ? 4'hd : _pms_pmx_T_84; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_86 = _T_108 ? 4'hc : _pms_pmx_T_85; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_87 = _T_107 ? 4'hb : _pms_pmx_T_86; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_88 = _T_106 ? 4'ha : _pms_pmx_T_87; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_89 = _T_105 ? 4'h9 : _pms_pmx_T_88; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_90 = _T_104 ? 4'h8 : _pms_pmx_T_89; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_91 = _T_103 ? 4'h7 : _pms_pmx_T_90; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_92 = _T_102 ? 4'h6 : _pms_pmx_T_91; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_93 = _T_101 ? 4'h5 : _pms_pmx_T_92; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_94 = _T_100 ? 4'h4 : _pms_pmx_T_93; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_95 = _T_99 ? 4'h3 : _pms_pmx_T_94; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_96 = _T_98 ? 4'h2 : _pms_pmx_T_95; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_97 = _T_97 ? 4'h1 : _pms_pmx_T_96; // @[Mux.scala 47:70]
  wire [3:0] pms_6 = _T_96 ? 4'h0 : _pms_pmx_T_97; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_98 = _T_126 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_99 = _T_125 ? 4'hd : _pms_pmx_T_98; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_100 = _T_124 ? 4'hc : _pms_pmx_T_99; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_101 = _T_123 ? 4'hb : _pms_pmx_T_100; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_102 = _T_122 ? 4'ha : _pms_pmx_T_101; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_103 = _T_121 ? 4'h9 : _pms_pmx_T_102; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_104 = _T_120 ? 4'h8 : _pms_pmx_T_103; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_105 = _T_119 ? 4'h7 : _pms_pmx_T_104; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_106 = _T_118 ? 4'h6 : _pms_pmx_T_105; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_107 = _T_117 ? 4'h5 : _pms_pmx_T_106; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_108 = _T_116 ? 4'h4 : _pms_pmx_T_107; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_109 = _T_115 ? 4'h3 : _pms_pmx_T_108; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_110 = _T_114 ? 4'h2 : _pms_pmx_T_109; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_111 = _T_113 ? 4'h1 : _pms_pmx_T_110; // @[Mux.scala 47:70]
  wire [3:0] pms_7 = _T_112 ? 4'h0 : _pms_pmx_T_111; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_112 = _T_142 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_113 = _T_141 ? 4'hd : _pms_pmx_T_112; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_114 = _T_140 ? 4'hc : _pms_pmx_T_113; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_115 = _T_139 ? 4'hb : _pms_pmx_T_114; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_116 = _T_138 ? 4'ha : _pms_pmx_T_115; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_117 = _T_137 ? 4'h9 : _pms_pmx_T_116; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_118 = _T_136 ? 4'h8 : _pms_pmx_T_117; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_119 = _T_135 ? 4'h7 : _pms_pmx_T_118; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_120 = _T_134 ? 4'h6 : _pms_pmx_T_119; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_121 = _T_133 ? 4'h5 : _pms_pmx_T_120; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_122 = _T_132 ? 4'h4 : _pms_pmx_T_121; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_123 = _T_131 ? 4'h3 : _pms_pmx_T_122; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_124 = _T_130 ? 4'h2 : _pms_pmx_T_123; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_125 = _T_129 ? 4'h1 : _pms_pmx_T_124; // @[Mux.scala 47:70]
  wire [3:0] pms_8 = _T_128 ? 4'h0 : _pms_pmx_T_125; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_126 = _T_158 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_127 = _T_157 ? 4'hd : _pms_pmx_T_126; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_128 = _T_156 ? 4'hc : _pms_pmx_T_127; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_129 = _T_155 ? 4'hb : _pms_pmx_T_128; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_130 = _T_154 ? 4'ha : _pms_pmx_T_129; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_131 = _T_153 ? 4'h9 : _pms_pmx_T_130; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_132 = _T_152 ? 4'h8 : _pms_pmx_T_131; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_133 = _T_151 ? 4'h7 : _pms_pmx_T_132; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_134 = _T_150 ? 4'h6 : _pms_pmx_T_133; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_135 = _T_149 ? 4'h5 : _pms_pmx_T_134; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_136 = _T_148 ? 4'h4 : _pms_pmx_T_135; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_137 = _T_147 ? 4'h3 : _pms_pmx_T_136; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_138 = _T_146 ? 4'h2 : _pms_pmx_T_137; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_139 = _T_145 ? 4'h1 : _pms_pmx_T_138; // @[Mux.scala 47:70]
  wire [3:0] pms_9 = _T_144 ? 4'h0 : _pms_pmx_T_139; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_140 = _T_174 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_141 = _T_173 ? 4'hd : _pms_pmx_T_140; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_142 = _T_172 ? 4'hc : _pms_pmx_T_141; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_143 = _T_171 ? 4'hb : _pms_pmx_T_142; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_144 = _T_170 ? 4'ha : _pms_pmx_T_143; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_145 = _T_169 ? 4'h9 : _pms_pmx_T_144; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_146 = _T_168 ? 4'h8 : _pms_pmx_T_145; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_147 = _T_167 ? 4'h7 : _pms_pmx_T_146; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_148 = _T_166 ? 4'h6 : _pms_pmx_T_147; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_149 = _T_165 ? 4'h5 : _pms_pmx_T_148; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_150 = _T_164 ? 4'h4 : _pms_pmx_T_149; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_151 = _T_163 ? 4'h3 : _pms_pmx_T_150; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_152 = _T_162 ? 4'h2 : _pms_pmx_T_151; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_153 = _T_161 ? 4'h1 : _pms_pmx_T_152; // @[Mux.scala 47:70]
  wire [3:0] pms_10 = _T_160 ? 4'h0 : _pms_pmx_T_153; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_154 = _T_190 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_155 = _T_189 ? 4'hd : _pms_pmx_T_154; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_156 = _T_188 ? 4'hc : _pms_pmx_T_155; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_157 = _T_187 ? 4'hb : _pms_pmx_T_156; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_158 = _T_186 ? 4'ha : _pms_pmx_T_157; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_159 = _T_185 ? 4'h9 : _pms_pmx_T_158; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_160 = _T_184 ? 4'h8 : _pms_pmx_T_159; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_161 = _T_183 ? 4'h7 : _pms_pmx_T_160; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_162 = _T_182 ? 4'h6 : _pms_pmx_T_161; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_163 = _T_181 ? 4'h5 : _pms_pmx_T_162; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_164 = _T_180 ? 4'h4 : _pms_pmx_T_163; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_165 = _T_179 ? 4'h3 : _pms_pmx_T_164; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_166 = _T_178 ? 4'h2 : _pms_pmx_T_165; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_167 = _T_177 ? 4'h1 : _pms_pmx_T_166; // @[Mux.scala 47:70]
  wire [3:0] pms_11 = _T_176 ? 4'h0 : _pms_pmx_T_167; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_168 = _T_206 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_169 = _T_205 ? 4'hd : _pms_pmx_T_168; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_170 = _T_204 ? 4'hc : _pms_pmx_T_169; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_171 = _T_203 ? 4'hb : _pms_pmx_T_170; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_172 = _T_202 ? 4'ha : _pms_pmx_T_171; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_173 = _T_201 ? 4'h9 : _pms_pmx_T_172; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_174 = _T_200 ? 4'h8 : _pms_pmx_T_173; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_175 = _T_199 ? 4'h7 : _pms_pmx_T_174; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_176 = _T_198 ? 4'h6 : _pms_pmx_T_175; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_177 = _T_197 ? 4'h5 : _pms_pmx_T_176; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_178 = _T_196 ? 4'h4 : _pms_pmx_T_177; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_179 = _T_195 ? 4'h3 : _pms_pmx_T_178; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_180 = _T_194 ? 4'h2 : _pms_pmx_T_179; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_181 = _T_193 ? 4'h1 : _pms_pmx_T_180; // @[Mux.scala 47:70]
  wire [3:0] pms_12 = _T_192 ? 4'h0 : _pms_pmx_T_181; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_182 = _T_222 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_183 = _T_221 ? 4'hd : _pms_pmx_T_182; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_184 = _T_220 ? 4'hc : _pms_pmx_T_183; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_185 = _T_219 ? 4'hb : _pms_pmx_T_184; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_186 = _T_218 ? 4'ha : _pms_pmx_T_185; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_187 = _T_217 ? 4'h9 : _pms_pmx_T_186; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_188 = _T_216 ? 4'h8 : _pms_pmx_T_187; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_189 = _T_215 ? 4'h7 : _pms_pmx_T_188; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_190 = _T_214 ? 4'h6 : _pms_pmx_T_189; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_191 = _T_213 ? 4'h5 : _pms_pmx_T_190; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_192 = _T_212 ? 4'h4 : _pms_pmx_T_191; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_193 = _T_211 ? 4'h3 : _pms_pmx_T_192; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_194 = _T_210 ? 4'h2 : _pms_pmx_T_193; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_195 = _T_209 ? 4'h1 : _pms_pmx_T_194; // @[Mux.scala 47:70]
  wire [3:0] pms_13 = _T_208 ? 4'h0 : _pms_pmx_T_195; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_196 = _T_238 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_197 = _T_237 ? 4'hd : _pms_pmx_T_196; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_198 = _T_236 ? 4'hc : _pms_pmx_T_197; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_199 = _T_235 ? 4'hb : _pms_pmx_T_198; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_200 = _T_234 ? 4'ha : _pms_pmx_T_199; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_201 = _T_233 ? 4'h9 : _pms_pmx_T_200; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_202 = _T_232 ? 4'h8 : _pms_pmx_T_201; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_203 = _T_231 ? 4'h7 : _pms_pmx_T_202; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_204 = _T_230 ? 4'h6 : _pms_pmx_T_203; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_205 = _T_229 ? 4'h5 : _pms_pmx_T_204; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_206 = _T_228 ? 4'h4 : _pms_pmx_T_205; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_207 = _T_227 ? 4'h3 : _pms_pmx_T_206; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_208 = _T_226 ? 4'h2 : _pms_pmx_T_207; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_209 = _T_225 ? 4'h1 : _pms_pmx_T_208; // @[Mux.scala 47:70]
  wire [3:0] pms_14 = _T_224 ? 4'h0 : _pms_pmx_T_209; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_210 = _T_254 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_211 = _T_253 ? 4'hd : _pms_pmx_T_210; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_212 = _T_252 ? 4'hc : _pms_pmx_T_211; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_213 = _T_251 ? 4'hb : _pms_pmx_T_212; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_214 = _T_250 ? 4'ha : _pms_pmx_T_213; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_215 = _T_249 ? 4'h9 : _pms_pmx_T_214; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_216 = _T_248 ? 4'h8 : _pms_pmx_T_215; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_217 = _T_247 ? 4'h7 : _pms_pmx_T_216; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_218 = _T_246 ? 4'h6 : _pms_pmx_T_217; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_219 = _T_245 ? 4'h5 : _pms_pmx_T_218; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_220 = _T_244 ? 4'h4 : _pms_pmx_T_219; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_221 = _T_243 ? 4'h3 : _pms_pmx_T_220; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_222 = _T_242 ? 4'h2 : _pms_pmx_T_221; // @[Mux.scala 47:70]
  wire [3:0] _pms_pmx_T_223 = _T_241 ? 4'h1 : _pms_pmx_T_222; // @[Mux.scala 47:70]
  wire [3:0] pms_15 = _T_240 ? 4'h0 : _pms_pmx_T_223; // @[Mux.scala 47:70]
  wire [31:0] _GEN_1 = 4'h1 == pms_0 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_2 = 4'h2 == pms_0 ? io_in_2_Im : _GEN_1; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_3 = 4'h3 == pms_0 ? io_in_3_Im : _GEN_2; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_4 = 4'h4 == pms_0 ? io_in_4_Im : _GEN_3; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_5 = 4'h5 == pms_0 ? io_in_5_Im : _GEN_4; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_6 = 4'h6 == pms_0 ? io_in_6_Im : _GEN_5; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_7 = 4'h7 == pms_0 ? io_in_7_Im : _GEN_6; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_8 = 4'h8 == pms_0 ? io_in_8_Im : _GEN_7; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_9 = 4'h9 == pms_0 ? io_in_9_Im : _GEN_8; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_10 = 4'ha == pms_0 ? io_in_10_Im : _GEN_9; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_11 = 4'hb == pms_0 ? io_in_11_Im : _GEN_10; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_12 = 4'hc == pms_0 ? io_in_12_Im : _GEN_11; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_13 = 4'hd == pms_0 ? io_in_13_Im : _GEN_12; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_14 = 4'he == pms_0 ? io_in_14_Im : _GEN_13; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_17 = 4'h1 == pms_0 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_18 = 4'h2 == pms_0 ? io_in_2_Re : _GEN_17; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_19 = 4'h3 == pms_0 ? io_in_3_Re : _GEN_18; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_20 = 4'h4 == pms_0 ? io_in_4_Re : _GEN_19; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_21 = 4'h5 == pms_0 ? io_in_5_Re : _GEN_20; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_22 = 4'h6 == pms_0 ? io_in_6_Re : _GEN_21; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_23 = 4'h7 == pms_0 ? io_in_7_Re : _GEN_22; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_24 = 4'h8 == pms_0 ? io_in_8_Re : _GEN_23; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_25 = 4'h9 == pms_0 ? io_in_9_Re : _GEN_24; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_26 = 4'ha == pms_0 ? io_in_10_Re : _GEN_25; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_27 = 4'hb == pms_0 ? io_in_11_Re : _GEN_26; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_28 = 4'hc == pms_0 ? io_in_12_Re : _GEN_27; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_29 = 4'hd == pms_0 ? io_in_13_Re : _GEN_28; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_30 = 4'he == pms_0 ? io_in_14_Re : _GEN_29; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_33 = 4'h1 == pms_1 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_34 = 4'h2 == pms_1 ? io_in_2_Im : _GEN_33; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_35 = 4'h3 == pms_1 ? io_in_3_Im : _GEN_34; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_36 = 4'h4 == pms_1 ? io_in_4_Im : _GEN_35; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_37 = 4'h5 == pms_1 ? io_in_5_Im : _GEN_36; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_38 = 4'h6 == pms_1 ? io_in_6_Im : _GEN_37; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_39 = 4'h7 == pms_1 ? io_in_7_Im : _GEN_38; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_40 = 4'h8 == pms_1 ? io_in_8_Im : _GEN_39; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_41 = 4'h9 == pms_1 ? io_in_9_Im : _GEN_40; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_42 = 4'ha == pms_1 ? io_in_10_Im : _GEN_41; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_43 = 4'hb == pms_1 ? io_in_11_Im : _GEN_42; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_44 = 4'hc == pms_1 ? io_in_12_Im : _GEN_43; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_45 = 4'hd == pms_1 ? io_in_13_Im : _GEN_44; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_46 = 4'he == pms_1 ? io_in_14_Im : _GEN_45; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_49 = 4'h1 == pms_1 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_50 = 4'h2 == pms_1 ? io_in_2_Re : _GEN_49; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_51 = 4'h3 == pms_1 ? io_in_3_Re : _GEN_50; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_52 = 4'h4 == pms_1 ? io_in_4_Re : _GEN_51; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_53 = 4'h5 == pms_1 ? io_in_5_Re : _GEN_52; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_54 = 4'h6 == pms_1 ? io_in_6_Re : _GEN_53; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_55 = 4'h7 == pms_1 ? io_in_7_Re : _GEN_54; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_56 = 4'h8 == pms_1 ? io_in_8_Re : _GEN_55; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_57 = 4'h9 == pms_1 ? io_in_9_Re : _GEN_56; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_58 = 4'ha == pms_1 ? io_in_10_Re : _GEN_57; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_59 = 4'hb == pms_1 ? io_in_11_Re : _GEN_58; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_60 = 4'hc == pms_1 ? io_in_12_Re : _GEN_59; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_61 = 4'hd == pms_1 ? io_in_13_Re : _GEN_60; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_62 = 4'he == pms_1 ? io_in_14_Re : _GEN_61; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_65 = 4'h1 == pms_2 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_66 = 4'h2 == pms_2 ? io_in_2_Im : _GEN_65; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_67 = 4'h3 == pms_2 ? io_in_3_Im : _GEN_66; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_68 = 4'h4 == pms_2 ? io_in_4_Im : _GEN_67; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_69 = 4'h5 == pms_2 ? io_in_5_Im : _GEN_68; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_70 = 4'h6 == pms_2 ? io_in_6_Im : _GEN_69; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_71 = 4'h7 == pms_2 ? io_in_7_Im : _GEN_70; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_72 = 4'h8 == pms_2 ? io_in_8_Im : _GEN_71; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_73 = 4'h9 == pms_2 ? io_in_9_Im : _GEN_72; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_74 = 4'ha == pms_2 ? io_in_10_Im : _GEN_73; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_75 = 4'hb == pms_2 ? io_in_11_Im : _GEN_74; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_76 = 4'hc == pms_2 ? io_in_12_Im : _GEN_75; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_77 = 4'hd == pms_2 ? io_in_13_Im : _GEN_76; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_78 = 4'he == pms_2 ? io_in_14_Im : _GEN_77; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_81 = 4'h1 == pms_2 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_82 = 4'h2 == pms_2 ? io_in_2_Re : _GEN_81; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_83 = 4'h3 == pms_2 ? io_in_3_Re : _GEN_82; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_84 = 4'h4 == pms_2 ? io_in_4_Re : _GEN_83; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_85 = 4'h5 == pms_2 ? io_in_5_Re : _GEN_84; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_86 = 4'h6 == pms_2 ? io_in_6_Re : _GEN_85; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_87 = 4'h7 == pms_2 ? io_in_7_Re : _GEN_86; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_88 = 4'h8 == pms_2 ? io_in_8_Re : _GEN_87; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_89 = 4'h9 == pms_2 ? io_in_9_Re : _GEN_88; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_90 = 4'ha == pms_2 ? io_in_10_Re : _GEN_89; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_91 = 4'hb == pms_2 ? io_in_11_Re : _GEN_90; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_92 = 4'hc == pms_2 ? io_in_12_Re : _GEN_91; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_93 = 4'hd == pms_2 ? io_in_13_Re : _GEN_92; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_94 = 4'he == pms_2 ? io_in_14_Re : _GEN_93; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_97 = 4'h1 == pms_3 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_98 = 4'h2 == pms_3 ? io_in_2_Im : _GEN_97; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_99 = 4'h3 == pms_3 ? io_in_3_Im : _GEN_98; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_100 = 4'h4 == pms_3 ? io_in_4_Im : _GEN_99; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_101 = 4'h5 == pms_3 ? io_in_5_Im : _GEN_100; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_102 = 4'h6 == pms_3 ? io_in_6_Im : _GEN_101; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_103 = 4'h7 == pms_3 ? io_in_7_Im : _GEN_102; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_104 = 4'h8 == pms_3 ? io_in_8_Im : _GEN_103; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_105 = 4'h9 == pms_3 ? io_in_9_Im : _GEN_104; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_106 = 4'ha == pms_3 ? io_in_10_Im : _GEN_105; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_107 = 4'hb == pms_3 ? io_in_11_Im : _GEN_106; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_108 = 4'hc == pms_3 ? io_in_12_Im : _GEN_107; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_109 = 4'hd == pms_3 ? io_in_13_Im : _GEN_108; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_110 = 4'he == pms_3 ? io_in_14_Im : _GEN_109; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_113 = 4'h1 == pms_3 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_114 = 4'h2 == pms_3 ? io_in_2_Re : _GEN_113; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_115 = 4'h3 == pms_3 ? io_in_3_Re : _GEN_114; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_116 = 4'h4 == pms_3 ? io_in_4_Re : _GEN_115; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_117 = 4'h5 == pms_3 ? io_in_5_Re : _GEN_116; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_118 = 4'h6 == pms_3 ? io_in_6_Re : _GEN_117; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_119 = 4'h7 == pms_3 ? io_in_7_Re : _GEN_118; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_120 = 4'h8 == pms_3 ? io_in_8_Re : _GEN_119; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_121 = 4'h9 == pms_3 ? io_in_9_Re : _GEN_120; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_122 = 4'ha == pms_3 ? io_in_10_Re : _GEN_121; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_123 = 4'hb == pms_3 ? io_in_11_Re : _GEN_122; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_124 = 4'hc == pms_3 ? io_in_12_Re : _GEN_123; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_125 = 4'hd == pms_3 ? io_in_13_Re : _GEN_124; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_126 = 4'he == pms_3 ? io_in_14_Re : _GEN_125; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_129 = 4'h1 == pms_4 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_130 = 4'h2 == pms_4 ? io_in_2_Im : _GEN_129; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_131 = 4'h3 == pms_4 ? io_in_3_Im : _GEN_130; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_132 = 4'h4 == pms_4 ? io_in_4_Im : _GEN_131; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_133 = 4'h5 == pms_4 ? io_in_5_Im : _GEN_132; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_134 = 4'h6 == pms_4 ? io_in_6_Im : _GEN_133; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_135 = 4'h7 == pms_4 ? io_in_7_Im : _GEN_134; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_136 = 4'h8 == pms_4 ? io_in_8_Im : _GEN_135; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_137 = 4'h9 == pms_4 ? io_in_9_Im : _GEN_136; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_138 = 4'ha == pms_4 ? io_in_10_Im : _GEN_137; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_139 = 4'hb == pms_4 ? io_in_11_Im : _GEN_138; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_140 = 4'hc == pms_4 ? io_in_12_Im : _GEN_139; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_141 = 4'hd == pms_4 ? io_in_13_Im : _GEN_140; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_142 = 4'he == pms_4 ? io_in_14_Im : _GEN_141; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_145 = 4'h1 == pms_4 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_146 = 4'h2 == pms_4 ? io_in_2_Re : _GEN_145; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_147 = 4'h3 == pms_4 ? io_in_3_Re : _GEN_146; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_148 = 4'h4 == pms_4 ? io_in_4_Re : _GEN_147; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_149 = 4'h5 == pms_4 ? io_in_5_Re : _GEN_148; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_150 = 4'h6 == pms_4 ? io_in_6_Re : _GEN_149; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_151 = 4'h7 == pms_4 ? io_in_7_Re : _GEN_150; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_152 = 4'h8 == pms_4 ? io_in_8_Re : _GEN_151; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_153 = 4'h9 == pms_4 ? io_in_9_Re : _GEN_152; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_154 = 4'ha == pms_4 ? io_in_10_Re : _GEN_153; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_155 = 4'hb == pms_4 ? io_in_11_Re : _GEN_154; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_156 = 4'hc == pms_4 ? io_in_12_Re : _GEN_155; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_157 = 4'hd == pms_4 ? io_in_13_Re : _GEN_156; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_158 = 4'he == pms_4 ? io_in_14_Re : _GEN_157; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_161 = 4'h1 == pms_5 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_162 = 4'h2 == pms_5 ? io_in_2_Im : _GEN_161; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_163 = 4'h3 == pms_5 ? io_in_3_Im : _GEN_162; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_164 = 4'h4 == pms_5 ? io_in_4_Im : _GEN_163; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_165 = 4'h5 == pms_5 ? io_in_5_Im : _GEN_164; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_166 = 4'h6 == pms_5 ? io_in_6_Im : _GEN_165; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_167 = 4'h7 == pms_5 ? io_in_7_Im : _GEN_166; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_168 = 4'h8 == pms_5 ? io_in_8_Im : _GEN_167; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_169 = 4'h9 == pms_5 ? io_in_9_Im : _GEN_168; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_170 = 4'ha == pms_5 ? io_in_10_Im : _GEN_169; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_171 = 4'hb == pms_5 ? io_in_11_Im : _GEN_170; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_172 = 4'hc == pms_5 ? io_in_12_Im : _GEN_171; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_173 = 4'hd == pms_5 ? io_in_13_Im : _GEN_172; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_174 = 4'he == pms_5 ? io_in_14_Im : _GEN_173; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_177 = 4'h1 == pms_5 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_178 = 4'h2 == pms_5 ? io_in_2_Re : _GEN_177; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_179 = 4'h3 == pms_5 ? io_in_3_Re : _GEN_178; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_180 = 4'h4 == pms_5 ? io_in_4_Re : _GEN_179; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_181 = 4'h5 == pms_5 ? io_in_5_Re : _GEN_180; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_182 = 4'h6 == pms_5 ? io_in_6_Re : _GEN_181; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_183 = 4'h7 == pms_5 ? io_in_7_Re : _GEN_182; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_184 = 4'h8 == pms_5 ? io_in_8_Re : _GEN_183; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_185 = 4'h9 == pms_5 ? io_in_9_Re : _GEN_184; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_186 = 4'ha == pms_5 ? io_in_10_Re : _GEN_185; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_187 = 4'hb == pms_5 ? io_in_11_Re : _GEN_186; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_188 = 4'hc == pms_5 ? io_in_12_Re : _GEN_187; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_189 = 4'hd == pms_5 ? io_in_13_Re : _GEN_188; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_190 = 4'he == pms_5 ? io_in_14_Re : _GEN_189; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_193 = 4'h1 == pms_6 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_194 = 4'h2 == pms_6 ? io_in_2_Im : _GEN_193; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_195 = 4'h3 == pms_6 ? io_in_3_Im : _GEN_194; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_196 = 4'h4 == pms_6 ? io_in_4_Im : _GEN_195; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_197 = 4'h5 == pms_6 ? io_in_5_Im : _GEN_196; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_198 = 4'h6 == pms_6 ? io_in_6_Im : _GEN_197; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_199 = 4'h7 == pms_6 ? io_in_7_Im : _GEN_198; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_200 = 4'h8 == pms_6 ? io_in_8_Im : _GEN_199; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_201 = 4'h9 == pms_6 ? io_in_9_Im : _GEN_200; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_202 = 4'ha == pms_6 ? io_in_10_Im : _GEN_201; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_203 = 4'hb == pms_6 ? io_in_11_Im : _GEN_202; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_204 = 4'hc == pms_6 ? io_in_12_Im : _GEN_203; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_205 = 4'hd == pms_6 ? io_in_13_Im : _GEN_204; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_206 = 4'he == pms_6 ? io_in_14_Im : _GEN_205; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_209 = 4'h1 == pms_6 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_210 = 4'h2 == pms_6 ? io_in_2_Re : _GEN_209; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_211 = 4'h3 == pms_6 ? io_in_3_Re : _GEN_210; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_212 = 4'h4 == pms_6 ? io_in_4_Re : _GEN_211; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_213 = 4'h5 == pms_6 ? io_in_5_Re : _GEN_212; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_214 = 4'h6 == pms_6 ? io_in_6_Re : _GEN_213; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_215 = 4'h7 == pms_6 ? io_in_7_Re : _GEN_214; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_216 = 4'h8 == pms_6 ? io_in_8_Re : _GEN_215; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_217 = 4'h9 == pms_6 ? io_in_9_Re : _GEN_216; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_218 = 4'ha == pms_6 ? io_in_10_Re : _GEN_217; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_219 = 4'hb == pms_6 ? io_in_11_Re : _GEN_218; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_220 = 4'hc == pms_6 ? io_in_12_Re : _GEN_219; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_221 = 4'hd == pms_6 ? io_in_13_Re : _GEN_220; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_222 = 4'he == pms_6 ? io_in_14_Re : _GEN_221; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_225 = 4'h1 == pms_7 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_226 = 4'h2 == pms_7 ? io_in_2_Im : _GEN_225; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_227 = 4'h3 == pms_7 ? io_in_3_Im : _GEN_226; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_228 = 4'h4 == pms_7 ? io_in_4_Im : _GEN_227; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_229 = 4'h5 == pms_7 ? io_in_5_Im : _GEN_228; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_230 = 4'h6 == pms_7 ? io_in_6_Im : _GEN_229; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_231 = 4'h7 == pms_7 ? io_in_7_Im : _GEN_230; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_232 = 4'h8 == pms_7 ? io_in_8_Im : _GEN_231; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_233 = 4'h9 == pms_7 ? io_in_9_Im : _GEN_232; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_234 = 4'ha == pms_7 ? io_in_10_Im : _GEN_233; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_235 = 4'hb == pms_7 ? io_in_11_Im : _GEN_234; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_236 = 4'hc == pms_7 ? io_in_12_Im : _GEN_235; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_237 = 4'hd == pms_7 ? io_in_13_Im : _GEN_236; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_238 = 4'he == pms_7 ? io_in_14_Im : _GEN_237; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_241 = 4'h1 == pms_7 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_242 = 4'h2 == pms_7 ? io_in_2_Re : _GEN_241; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_243 = 4'h3 == pms_7 ? io_in_3_Re : _GEN_242; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_244 = 4'h4 == pms_7 ? io_in_4_Re : _GEN_243; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_245 = 4'h5 == pms_7 ? io_in_5_Re : _GEN_244; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_246 = 4'h6 == pms_7 ? io_in_6_Re : _GEN_245; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_247 = 4'h7 == pms_7 ? io_in_7_Re : _GEN_246; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_248 = 4'h8 == pms_7 ? io_in_8_Re : _GEN_247; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_249 = 4'h9 == pms_7 ? io_in_9_Re : _GEN_248; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_250 = 4'ha == pms_7 ? io_in_10_Re : _GEN_249; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_251 = 4'hb == pms_7 ? io_in_11_Re : _GEN_250; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_252 = 4'hc == pms_7 ? io_in_12_Re : _GEN_251; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_253 = 4'hd == pms_7 ? io_in_13_Re : _GEN_252; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_254 = 4'he == pms_7 ? io_in_14_Re : _GEN_253; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_257 = 4'h1 == pms_8 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_258 = 4'h2 == pms_8 ? io_in_2_Im : _GEN_257; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_259 = 4'h3 == pms_8 ? io_in_3_Im : _GEN_258; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_260 = 4'h4 == pms_8 ? io_in_4_Im : _GEN_259; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_261 = 4'h5 == pms_8 ? io_in_5_Im : _GEN_260; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_262 = 4'h6 == pms_8 ? io_in_6_Im : _GEN_261; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_263 = 4'h7 == pms_8 ? io_in_7_Im : _GEN_262; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_264 = 4'h8 == pms_8 ? io_in_8_Im : _GEN_263; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_265 = 4'h9 == pms_8 ? io_in_9_Im : _GEN_264; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_266 = 4'ha == pms_8 ? io_in_10_Im : _GEN_265; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_267 = 4'hb == pms_8 ? io_in_11_Im : _GEN_266; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_268 = 4'hc == pms_8 ? io_in_12_Im : _GEN_267; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_269 = 4'hd == pms_8 ? io_in_13_Im : _GEN_268; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_270 = 4'he == pms_8 ? io_in_14_Im : _GEN_269; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_273 = 4'h1 == pms_8 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_274 = 4'h2 == pms_8 ? io_in_2_Re : _GEN_273; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_275 = 4'h3 == pms_8 ? io_in_3_Re : _GEN_274; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_276 = 4'h4 == pms_8 ? io_in_4_Re : _GEN_275; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_277 = 4'h5 == pms_8 ? io_in_5_Re : _GEN_276; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_278 = 4'h6 == pms_8 ? io_in_6_Re : _GEN_277; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_279 = 4'h7 == pms_8 ? io_in_7_Re : _GEN_278; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_280 = 4'h8 == pms_8 ? io_in_8_Re : _GEN_279; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_281 = 4'h9 == pms_8 ? io_in_9_Re : _GEN_280; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_282 = 4'ha == pms_8 ? io_in_10_Re : _GEN_281; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_283 = 4'hb == pms_8 ? io_in_11_Re : _GEN_282; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_284 = 4'hc == pms_8 ? io_in_12_Re : _GEN_283; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_285 = 4'hd == pms_8 ? io_in_13_Re : _GEN_284; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_286 = 4'he == pms_8 ? io_in_14_Re : _GEN_285; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_289 = 4'h1 == pms_9 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_290 = 4'h2 == pms_9 ? io_in_2_Im : _GEN_289; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_291 = 4'h3 == pms_9 ? io_in_3_Im : _GEN_290; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_292 = 4'h4 == pms_9 ? io_in_4_Im : _GEN_291; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_293 = 4'h5 == pms_9 ? io_in_5_Im : _GEN_292; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_294 = 4'h6 == pms_9 ? io_in_6_Im : _GEN_293; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_295 = 4'h7 == pms_9 ? io_in_7_Im : _GEN_294; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_296 = 4'h8 == pms_9 ? io_in_8_Im : _GEN_295; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_297 = 4'h9 == pms_9 ? io_in_9_Im : _GEN_296; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_298 = 4'ha == pms_9 ? io_in_10_Im : _GEN_297; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_299 = 4'hb == pms_9 ? io_in_11_Im : _GEN_298; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_300 = 4'hc == pms_9 ? io_in_12_Im : _GEN_299; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_301 = 4'hd == pms_9 ? io_in_13_Im : _GEN_300; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_302 = 4'he == pms_9 ? io_in_14_Im : _GEN_301; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_305 = 4'h1 == pms_9 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_306 = 4'h2 == pms_9 ? io_in_2_Re : _GEN_305; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_307 = 4'h3 == pms_9 ? io_in_3_Re : _GEN_306; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_308 = 4'h4 == pms_9 ? io_in_4_Re : _GEN_307; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_309 = 4'h5 == pms_9 ? io_in_5_Re : _GEN_308; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_310 = 4'h6 == pms_9 ? io_in_6_Re : _GEN_309; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_311 = 4'h7 == pms_9 ? io_in_7_Re : _GEN_310; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_312 = 4'h8 == pms_9 ? io_in_8_Re : _GEN_311; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_313 = 4'h9 == pms_9 ? io_in_9_Re : _GEN_312; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_314 = 4'ha == pms_9 ? io_in_10_Re : _GEN_313; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_315 = 4'hb == pms_9 ? io_in_11_Re : _GEN_314; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_316 = 4'hc == pms_9 ? io_in_12_Re : _GEN_315; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_317 = 4'hd == pms_9 ? io_in_13_Re : _GEN_316; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_318 = 4'he == pms_9 ? io_in_14_Re : _GEN_317; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_321 = 4'h1 == pms_10 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_322 = 4'h2 == pms_10 ? io_in_2_Im : _GEN_321; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_323 = 4'h3 == pms_10 ? io_in_3_Im : _GEN_322; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_324 = 4'h4 == pms_10 ? io_in_4_Im : _GEN_323; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_325 = 4'h5 == pms_10 ? io_in_5_Im : _GEN_324; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_326 = 4'h6 == pms_10 ? io_in_6_Im : _GEN_325; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_327 = 4'h7 == pms_10 ? io_in_7_Im : _GEN_326; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_328 = 4'h8 == pms_10 ? io_in_8_Im : _GEN_327; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_329 = 4'h9 == pms_10 ? io_in_9_Im : _GEN_328; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_330 = 4'ha == pms_10 ? io_in_10_Im : _GEN_329; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_331 = 4'hb == pms_10 ? io_in_11_Im : _GEN_330; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_332 = 4'hc == pms_10 ? io_in_12_Im : _GEN_331; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_333 = 4'hd == pms_10 ? io_in_13_Im : _GEN_332; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_334 = 4'he == pms_10 ? io_in_14_Im : _GEN_333; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_337 = 4'h1 == pms_10 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_338 = 4'h2 == pms_10 ? io_in_2_Re : _GEN_337; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_339 = 4'h3 == pms_10 ? io_in_3_Re : _GEN_338; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_340 = 4'h4 == pms_10 ? io_in_4_Re : _GEN_339; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_341 = 4'h5 == pms_10 ? io_in_5_Re : _GEN_340; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_342 = 4'h6 == pms_10 ? io_in_6_Re : _GEN_341; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_343 = 4'h7 == pms_10 ? io_in_7_Re : _GEN_342; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_344 = 4'h8 == pms_10 ? io_in_8_Re : _GEN_343; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_345 = 4'h9 == pms_10 ? io_in_9_Re : _GEN_344; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_346 = 4'ha == pms_10 ? io_in_10_Re : _GEN_345; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_347 = 4'hb == pms_10 ? io_in_11_Re : _GEN_346; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_348 = 4'hc == pms_10 ? io_in_12_Re : _GEN_347; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_349 = 4'hd == pms_10 ? io_in_13_Re : _GEN_348; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_350 = 4'he == pms_10 ? io_in_14_Re : _GEN_349; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_353 = 4'h1 == pms_11 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_354 = 4'h2 == pms_11 ? io_in_2_Im : _GEN_353; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_355 = 4'h3 == pms_11 ? io_in_3_Im : _GEN_354; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_356 = 4'h4 == pms_11 ? io_in_4_Im : _GEN_355; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_357 = 4'h5 == pms_11 ? io_in_5_Im : _GEN_356; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_358 = 4'h6 == pms_11 ? io_in_6_Im : _GEN_357; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_359 = 4'h7 == pms_11 ? io_in_7_Im : _GEN_358; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_360 = 4'h8 == pms_11 ? io_in_8_Im : _GEN_359; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_361 = 4'h9 == pms_11 ? io_in_9_Im : _GEN_360; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_362 = 4'ha == pms_11 ? io_in_10_Im : _GEN_361; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_363 = 4'hb == pms_11 ? io_in_11_Im : _GEN_362; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_364 = 4'hc == pms_11 ? io_in_12_Im : _GEN_363; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_365 = 4'hd == pms_11 ? io_in_13_Im : _GEN_364; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_366 = 4'he == pms_11 ? io_in_14_Im : _GEN_365; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_369 = 4'h1 == pms_11 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_370 = 4'h2 == pms_11 ? io_in_2_Re : _GEN_369; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_371 = 4'h3 == pms_11 ? io_in_3_Re : _GEN_370; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_372 = 4'h4 == pms_11 ? io_in_4_Re : _GEN_371; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_373 = 4'h5 == pms_11 ? io_in_5_Re : _GEN_372; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_374 = 4'h6 == pms_11 ? io_in_6_Re : _GEN_373; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_375 = 4'h7 == pms_11 ? io_in_7_Re : _GEN_374; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_376 = 4'h8 == pms_11 ? io_in_8_Re : _GEN_375; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_377 = 4'h9 == pms_11 ? io_in_9_Re : _GEN_376; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_378 = 4'ha == pms_11 ? io_in_10_Re : _GEN_377; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_379 = 4'hb == pms_11 ? io_in_11_Re : _GEN_378; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_380 = 4'hc == pms_11 ? io_in_12_Re : _GEN_379; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_381 = 4'hd == pms_11 ? io_in_13_Re : _GEN_380; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_382 = 4'he == pms_11 ? io_in_14_Re : _GEN_381; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_385 = 4'h1 == pms_12 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_386 = 4'h2 == pms_12 ? io_in_2_Im : _GEN_385; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_387 = 4'h3 == pms_12 ? io_in_3_Im : _GEN_386; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_388 = 4'h4 == pms_12 ? io_in_4_Im : _GEN_387; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_389 = 4'h5 == pms_12 ? io_in_5_Im : _GEN_388; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_390 = 4'h6 == pms_12 ? io_in_6_Im : _GEN_389; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_391 = 4'h7 == pms_12 ? io_in_7_Im : _GEN_390; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_392 = 4'h8 == pms_12 ? io_in_8_Im : _GEN_391; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_393 = 4'h9 == pms_12 ? io_in_9_Im : _GEN_392; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_394 = 4'ha == pms_12 ? io_in_10_Im : _GEN_393; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_395 = 4'hb == pms_12 ? io_in_11_Im : _GEN_394; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_396 = 4'hc == pms_12 ? io_in_12_Im : _GEN_395; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_397 = 4'hd == pms_12 ? io_in_13_Im : _GEN_396; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_398 = 4'he == pms_12 ? io_in_14_Im : _GEN_397; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_401 = 4'h1 == pms_12 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_402 = 4'h2 == pms_12 ? io_in_2_Re : _GEN_401; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_403 = 4'h3 == pms_12 ? io_in_3_Re : _GEN_402; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_404 = 4'h4 == pms_12 ? io_in_4_Re : _GEN_403; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_405 = 4'h5 == pms_12 ? io_in_5_Re : _GEN_404; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_406 = 4'h6 == pms_12 ? io_in_6_Re : _GEN_405; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_407 = 4'h7 == pms_12 ? io_in_7_Re : _GEN_406; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_408 = 4'h8 == pms_12 ? io_in_8_Re : _GEN_407; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_409 = 4'h9 == pms_12 ? io_in_9_Re : _GEN_408; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_410 = 4'ha == pms_12 ? io_in_10_Re : _GEN_409; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_411 = 4'hb == pms_12 ? io_in_11_Re : _GEN_410; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_412 = 4'hc == pms_12 ? io_in_12_Re : _GEN_411; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_413 = 4'hd == pms_12 ? io_in_13_Re : _GEN_412; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_414 = 4'he == pms_12 ? io_in_14_Re : _GEN_413; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_417 = 4'h1 == pms_13 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_418 = 4'h2 == pms_13 ? io_in_2_Im : _GEN_417; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_419 = 4'h3 == pms_13 ? io_in_3_Im : _GEN_418; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_420 = 4'h4 == pms_13 ? io_in_4_Im : _GEN_419; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_421 = 4'h5 == pms_13 ? io_in_5_Im : _GEN_420; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_422 = 4'h6 == pms_13 ? io_in_6_Im : _GEN_421; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_423 = 4'h7 == pms_13 ? io_in_7_Im : _GEN_422; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_424 = 4'h8 == pms_13 ? io_in_8_Im : _GEN_423; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_425 = 4'h9 == pms_13 ? io_in_9_Im : _GEN_424; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_426 = 4'ha == pms_13 ? io_in_10_Im : _GEN_425; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_427 = 4'hb == pms_13 ? io_in_11_Im : _GEN_426; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_428 = 4'hc == pms_13 ? io_in_12_Im : _GEN_427; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_429 = 4'hd == pms_13 ? io_in_13_Im : _GEN_428; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_430 = 4'he == pms_13 ? io_in_14_Im : _GEN_429; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_433 = 4'h1 == pms_13 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_434 = 4'h2 == pms_13 ? io_in_2_Re : _GEN_433; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_435 = 4'h3 == pms_13 ? io_in_3_Re : _GEN_434; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_436 = 4'h4 == pms_13 ? io_in_4_Re : _GEN_435; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_437 = 4'h5 == pms_13 ? io_in_5_Re : _GEN_436; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_438 = 4'h6 == pms_13 ? io_in_6_Re : _GEN_437; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_439 = 4'h7 == pms_13 ? io_in_7_Re : _GEN_438; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_440 = 4'h8 == pms_13 ? io_in_8_Re : _GEN_439; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_441 = 4'h9 == pms_13 ? io_in_9_Re : _GEN_440; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_442 = 4'ha == pms_13 ? io_in_10_Re : _GEN_441; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_443 = 4'hb == pms_13 ? io_in_11_Re : _GEN_442; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_444 = 4'hc == pms_13 ? io_in_12_Re : _GEN_443; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_445 = 4'hd == pms_13 ? io_in_13_Re : _GEN_444; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_446 = 4'he == pms_13 ? io_in_14_Re : _GEN_445; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_449 = 4'h1 == pms_14 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_450 = 4'h2 == pms_14 ? io_in_2_Im : _GEN_449; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_451 = 4'h3 == pms_14 ? io_in_3_Im : _GEN_450; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_452 = 4'h4 == pms_14 ? io_in_4_Im : _GEN_451; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_453 = 4'h5 == pms_14 ? io_in_5_Im : _GEN_452; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_454 = 4'h6 == pms_14 ? io_in_6_Im : _GEN_453; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_455 = 4'h7 == pms_14 ? io_in_7_Im : _GEN_454; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_456 = 4'h8 == pms_14 ? io_in_8_Im : _GEN_455; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_457 = 4'h9 == pms_14 ? io_in_9_Im : _GEN_456; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_458 = 4'ha == pms_14 ? io_in_10_Im : _GEN_457; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_459 = 4'hb == pms_14 ? io_in_11_Im : _GEN_458; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_460 = 4'hc == pms_14 ? io_in_12_Im : _GEN_459; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_461 = 4'hd == pms_14 ? io_in_13_Im : _GEN_460; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_462 = 4'he == pms_14 ? io_in_14_Im : _GEN_461; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_465 = 4'h1 == pms_14 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_466 = 4'h2 == pms_14 ? io_in_2_Re : _GEN_465; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_467 = 4'h3 == pms_14 ? io_in_3_Re : _GEN_466; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_468 = 4'h4 == pms_14 ? io_in_4_Re : _GEN_467; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_469 = 4'h5 == pms_14 ? io_in_5_Re : _GEN_468; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_470 = 4'h6 == pms_14 ? io_in_6_Re : _GEN_469; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_471 = 4'h7 == pms_14 ? io_in_7_Re : _GEN_470; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_472 = 4'h8 == pms_14 ? io_in_8_Re : _GEN_471; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_473 = 4'h9 == pms_14 ? io_in_9_Re : _GEN_472; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_474 = 4'ha == pms_14 ? io_in_10_Re : _GEN_473; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_475 = 4'hb == pms_14 ? io_in_11_Re : _GEN_474; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_476 = 4'hc == pms_14 ? io_in_12_Re : _GEN_475; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_477 = 4'hd == pms_14 ? io_in_13_Re : _GEN_476; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_478 = 4'he == pms_14 ? io_in_14_Re : _GEN_477; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_481 = 4'h1 == pms_15 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_482 = 4'h2 == pms_15 ? io_in_2_Im : _GEN_481; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_483 = 4'h3 == pms_15 ? io_in_3_Im : _GEN_482; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_484 = 4'h4 == pms_15 ? io_in_4_Im : _GEN_483; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_485 = 4'h5 == pms_15 ? io_in_5_Im : _GEN_484; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_486 = 4'h6 == pms_15 ? io_in_6_Im : _GEN_485; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_487 = 4'h7 == pms_15 ? io_in_7_Im : _GEN_486; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_488 = 4'h8 == pms_15 ? io_in_8_Im : _GEN_487; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_489 = 4'h9 == pms_15 ? io_in_9_Im : _GEN_488; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_490 = 4'ha == pms_15 ? io_in_10_Im : _GEN_489; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_491 = 4'hb == pms_15 ? io_in_11_Im : _GEN_490; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_492 = 4'hc == pms_15 ? io_in_12_Im : _GEN_491; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_493 = 4'hd == pms_15 ? io_in_13_Im : _GEN_492; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_494 = 4'he == pms_15 ? io_in_14_Im : _GEN_493; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_497 = 4'h1 == pms_15 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_498 = 4'h2 == pms_15 ? io_in_2_Re : _GEN_497; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_499 = 4'h3 == pms_15 ? io_in_3_Re : _GEN_498; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_500 = 4'h4 == pms_15 ? io_in_4_Re : _GEN_499; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_501 = 4'h5 == pms_15 ? io_in_5_Re : _GEN_500; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_502 = 4'h6 == pms_15 ? io_in_6_Re : _GEN_501; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_503 = 4'h7 == pms_15 ? io_in_7_Re : _GEN_502; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_504 = 4'h8 == pms_15 ? io_in_8_Re : _GEN_503; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_505 = 4'h9 == pms_15 ? io_in_9_Re : _GEN_504; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_506 = 4'ha == pms_15 ? io_in_10_Re : _GEN_505; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_507 = 4'hb == pms_15 ? io_in_11_Re : _GEN_506; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_508 = 4'hc == pms_15 ? io_in_12_Re : _GEN_507; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_509 = 4'hd == pms_15 ? io_in_13_Re : _GEN_508; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_510 = 4'he == pms_15 ? io_in_14_Re : _GEN_509; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_0_Re = 4'hf == pms_0 ? io_in_15_Re : _GEN_30; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_0_Im = 4'hf == pms_0 ? io_in_15_Im : _GEN_14; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_1_Re = 4'hf == pms_1 ? io_in_15_Re : _GEN_62; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_1_Im = 4'hf == pms_1 ? io_in_15_Im : _GEN_46; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_2_Re = 4'hf == pms_2 ? io_in_15_Re : _GEN_94; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_2_Im = 4'hf == pms_2 ? io_in_15_Im : _GEN_78; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_3_Re = 4'hf == pms_3 ? io_in_15_Re : _GEN_126; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_3_Im = 4'hf == pms_3 ? io_in_15_Im : _GEN_110; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_4_Re = 4'hf == pms_4 ? io_in_15_Re : _GEN_158; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_4_Im = 4'hf == pms_4 ? io_in_15_Im : _GEN_142; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_5_Re = 4'hf == pms_5 ? io_in_15_Re : _GEN_190; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_5_Im = 4'hf == pms_5 ? io_in_15_Im : _GEN_174; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_6_Re = 4'hf == pms_6 ? io_in_15_Re : _GEN_222; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_6_Im = 4'hf == pms_6 ? io_in_15_Im : _GEN_206; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_7_Re = 4'hf == pms_7 ? io_in_15_Re : _GEN_254; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_7_Im = 4'hf == pms_7 ? io_in_15_Im : _GEN_238; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_8_Re = 4'hf == pms_8 ? io_in_15_Re : _GEN_286; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_8_Im = 4'hf == pms_8 ? io_in_15_Im : _GEN_270; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_9_Re = 4'hf == pms_9 ? io_in_15_Re : _GEN_318; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_9_Im = 4'hf == pms_9 ? io_in_15_Im : _GEN_302; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_10_Re = 4'hf == pms_10 ? io_in_15_Re : _GEN_350; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_10_Im = 4'hf == pms_10 ? io_in_15_Im : _GEN_334; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_11_Re = 4'hf == pms_11 ? io_in_15_Re : _GEN_382; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_11_Im = 4'hf == pms_11 ? io_in_15_Im : _GEN_366; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_12_Re = 4'hf == pms_12 ? io_in_15_Re : _GEN_414; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_12_Im = 4'hf == pms_12 ? io_in_15_Im : _GEN_398; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_13_Re = 4'hf == pms_13 ? io_in_15_Re : _GEN_446; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_13_Im = 4'hf == pms_13 ? io_in_15_Im : _GEN_430; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_14_Re = 4'hf == pms_14 ? io_in_15_Re : _GEN_478; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_14_Im = 4'hf == pms_14 ? io_in_15_Im : _GEN_462; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_15_Re = 4'hf == pms_15 ? io_in_15_Re : _GEN_510; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_15_Im = 4'hf == pms_15 ? io_in_15_Im : _GEN_494; // @[FFTDesigns.scala 3203:{17,17}]
endmodule
module M0_Config_ROM(
  input        io_in_cnt,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2,
  output [1:0] io_out_3,
  output [1:0] io_out_4,
  output [1:0] io_out_5,
  output [1:0] io_out_6,
  output [1:0] io_out_7,
  output [1:0] io_out_8,
  output [1:0] io_out_9,
  output [1:0] io_out_10,
  output [1:0] io_out_11,
  output [1:0] io_out_12,
  output [1:0] io_out_13,
  output [1:0] io_out_14,
  output [1:0] io_out_15
);
  assign io_out_0 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_1 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_2 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_3 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_4 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_5 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_6 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_7 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_8 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_9 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_10 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_11 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_12 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_13 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_14 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_15 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3227:{17,17}]
endmodule
module M1_Config_ROM(
  input        io_in_cnt,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2,
  output [1:0] io_out_3,
  output [1:0] io_out_4,
  output [1:0] io_out_5,
  output [1:0] io_out_6,
  output [1:0] io_out_7,
  output [1:0] io_out_8,
  output [1:0] io_out_9,
  output [1:0] io_out_10,
  output [1:0] io_out_11,
  output [1:0] io_out_12,
  output [1:0] io_out_13,
  output [1:0] io_out_14,
  output [1:0] io_out_15
);
  assign io_out_0 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_1 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_2 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_3 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_4 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_5 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_6 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_7 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_8 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_9 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_10 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_11 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_12 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_13 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_14 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_15 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
endmodule
module Streaming_Permute_Config(
  input        io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11,
  output [3:0] io_out_12,
  output [3:0] io_out_13,
  output [3:0] io_out_14
);
  assign io_out_0 = io_in_cnt ? 4'h1 : 4'h0; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_1 = io_in_cnt ? 4'h0 : 4'h1; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_2 = io_in_cnt ? 4'h9 : 4'h8; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_3 = io_in_cnt ? 4'h8 : 4'h9; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_4 = io_in_cnt ? 4'h5 : 4'h4; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_5 = io_in_cnt ? 4'h4 : 4'h5; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_6 = io_in_cnt ? 4'hd : 4'hc; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_7 = io_in_cnt ? 4'hc : 4'hd; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_8 = io_in_cnt ? 4'h3 : 4'h2; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_9 = io_in_cnt ? 4'h2 : 4'h3; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_10 = io_in_cnt ? 4'hb : 4'ha; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_11 = io_in_cnt ? 4'ha : 4'hb; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_12 = io_in_cnt ? 4'h7 : 4'h6; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_13 = io_in_cnt ? 4'h6 : 4'h7; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_14 = io_in_cnt ? 4'hf : 4'he; // @[FFTDesigns.scala 3273:{17,17}]
endmodule
module PermutationsWithStreaming(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_16_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_16_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_16_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_17_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_17_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_18_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_18_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_19_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_19_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_20_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_20_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_21_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_21_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_22_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_22_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_23_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_23_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_24_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_24_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_25_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_25_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_26_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_26_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_27_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_27_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_28_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_28_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_29_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_29_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_30_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_30_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_31_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_31_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_8_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_8_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_9_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_9_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_10_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_10_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_11_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_11_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_12_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_12_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_13_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_13_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_14_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_14_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_15_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_15_Im; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_7; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_8; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_9; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_10; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_11; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_12; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_13; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_14; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2641:26]
  wire  M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_8; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_9; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_10; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_11; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_12; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_13; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_14; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_15; // @[FFTDesigns.scala 2642:27]
  wire  M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_8; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_9; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_10; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_11; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_12; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_13; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_14; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_15; // @[FFTDesigns.scala 2643:27]
  wire  Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2644:29]
  reg  offset_switch; // @[FFTDesigns.scala 2627:28]
  wire [4:0] _T = {io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2628:19]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2628:26]
  reg  cnt; // @[FFTDesigns.scala 2645:22]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2649:26]
  wire  _GEN_1 = cnt ? 1'h0 : cnt + 1'h1; // @[FFTDesigns.scala 2647:32 2648:13 2651:13]
  wire  _GEN_2 = cnt ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2647:32 2649:23 2652:23]
  wire [2:0] _T_6 = 2'h2 * _offset_switch_T; // @[FFTDesigns.scala 2661:54]
  wire [2:0] _GEN_214 = {{1'd0}, M0_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_8 = _GEN_214 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_9 = 2'h2 * offset_switch; // @[FFTDesigns.scala 2662:41]
  wire [2:0] _GEN_215 = {{2'd0}, cnt}; // @[FFTDesigns.scala 2662:31]
  wire [2:0] _T_11 = _GEN_215 + _T_9; // @[FFTDesigns.scala 2662:31]
  wire [2:0] _T_15 = _GEN_215 + _T_6; // @[FFTDesigns.scala 2664:31]
  wire [2:0] _GEN_217 = {{1'd0}, M1_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_18 = _GEN_217 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_218 = {{1'd0}, M0_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_22 = _GEN_218 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_221 = {{1'd0}, M1_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_32 = _GEN_221 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_222 = {{1'd0}, M0_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_36 = _GEN_222 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_225 = {{1'd0}, M1_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_46 = _GEN_225 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_226 = {{1'd0}, M0_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_50 = _GEN_226 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_229 = {{1'd0}, M1_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_60 = _GEN_229 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_230 = {{1'd0}, M0_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_64 = _GEN_230 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_233 = {{1'd0}, M1_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_74 = _GEN_233 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_234 = {{1'd0}, M0_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_78 = _GEN_234 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_237 = {{1'd0}, M1_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_88 = _GEN_237 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_238 = {{1'd0}, M0_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_92 = _GEN_238 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_241 = {{1'd0}, M1_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_102 = _GEN_241 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_242 = {{1'd0}, M0_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_106 = _GEN_242 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_245 = {{1'd0}, M1_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_116 = _GEN_245 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_246 = {{1'd0}, M0_Config_ROM_io_out_8}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_120 = _GEN_246 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_249 = {{1'd0}, M1_Config_ROM_io_out_8}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_130 = _GEN_249 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_250 = {{1'd0}, M0_Config_ROM_io_out_9}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_134 = _GEN_250 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_253 = {{1'd0}, M1_Config_ROM_io_out_9}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_144 = _GEN_253 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_254 = {{1'd0}, M0_Config_ROM_io_out_10}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_148 = _GEN_254 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_257 = {{1'd0}, M1_Config_ROM_io_out_10}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_158 = _GEN_257 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_258 = {{1'd0}, M0_Config_ROM_io_out_11}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_162 = _GEN_258 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_261 = {{1'd0}, M1_Config_ROM_io_out_11}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_172 = _GEN_261 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_262 = {{1'd0}, M0_Config_ROM_io_out_12}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_176 = _GEN_262 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_265 = {{1'd0}, M1_Config_ROM_io_out_12}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_186 = _GEN_265 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_266 = {{1'd0}, M0_Config_ROM_io_out_13}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_190 = _GEN_266 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_269 = {{1'd0}, M1_Config_ROM_io_out_13}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_200 = _GEN_269 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_270 = {{1'd0}, M0_Config_ROM_io_out_14}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_204 = _GEN_270 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_273 = {{1'd0}, M1_Config_ROM_io_out_14}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_214 = _GEN_273 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_274 = {{1'd0}, M0_Config_ROM_io_out_15}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_218 = _GEN_274 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_277 = {{1'd0}, M1_Config_ROM_io_out_15}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_228 = _GEN_277 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire  _GEN_3 = _T_1 & _GEN_1; // @[FFTDesigns.scala 2646:30 2692:11]
  wire [2:0] _GEN_6 = _T_1 ? _T_8 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_7 = _T_1 ? _T_11 : 3'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  wire [2:0] _GEN_10 = _T_1 ? _T_15 : 3'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  wire [2:0] _GEN_11 = _T_1 ? _T_18 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_19 = _T_1 ? _T_22 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_24 = _T_1 ? _T_32 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_32 = _T_1 ? _T_36 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_37 = _T_1 ? _T_46 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_45 = _T_1 ? _T_50 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_50 = _T_1 ? _T_60 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_58 = _T_1 ? _T_64 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_63 = _T_1 ? _T_74 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_71 = _T_1 ? _T_78 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_76 = _T_1 ? _T_88 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_84 = _T_1 ? _T_92 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_89 = _T_1 ? _T_102 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_97 = _T_1 ? _T_106 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_102 = _T_1 ? _T_116 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_110 = _T_1 ? _T_120 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_115 = _T_1 ? _T_130 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_123 = _T_1 ? _T_134 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_128 = _T_1 ? _T_144 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_136 = _T_1 ? _T_148 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_141 = _T_1 ? _T_158 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_149 = _T_1 ? _T_162 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_154 = _T_1 ? _T_172 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_162 = _T_1 ? _T_176 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_167 = _T_1 ? _T_186 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_175 = _T_1 ? _T_190 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_180 = _T_1 ? _T_200 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_188 = _T_1 ? _T_204 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_193 = _T_1 ? _T_214 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_201 = _T_1 ? _T_218 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_206 = _T_1 ? _T_228 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  RAM_Block RAM_Block ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block RAM_Block_1 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block RAM_Block_2 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block RAM_Block_3 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block RAM_Block_4 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block RAM_Block_5 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block RAM_Block_6 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block RAM_Block_7 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block RAM_Block_8 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block RAM_Block_9 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block RAM_Block_10 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block RAM_Block_11 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block RAM_Block_12 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block RAM_Block_13 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block RAM_Block_14 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block RAM_Block_15 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  RAM_Block RAM_Block_16 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_16_clock),
    .io_in_raddr(RAM_Block_16_io_in_raddr),
    .io_in_waddr(RAM_Block_16_io_in_waddr),
    .io_in_data_Re(RAM_Block_16_io_in_data_Re),
    .io_in_data_Im(RAM_Block_16_io_in_data_Im),
    .io_re(RAM_Block_16_io_re),
    .io_wr(RAM_Block_16_io_wr),
    .io_en(RAM_Block_16_io_en),
    .io_out_data_Re(RAM_Block_16_io_out_data_Re),
    .io_out_data_Im(RAM_Block_16_io_out_data_Im)
  );
  RAM_Block RAM_Block_17 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_17_clock),
    .io_in_raddr(RAM_Block_17_io_in_raddr),
    .io_in_waddr(RAM_Block_17_io_in_waddr),
    .io_in_data_Re(RAM_Block_17_io_in_data_Re),
    .io_in_data_Im(RAM_Block_17_io_in_data_Im),
    .io_re(RAM_Block_17_io_re),
    .io_wr(RAM_Block_17_io_wr),
    .io_en(RAM_Block_17_io_en),
    .io_out_data_Re(RAM_Block_17_io_out_data_Re),
    .io_out_data_Im(RAM_Block_17_io_out_data_Im)
  );
  RAM_Block RAM_Block_18 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_18_clock),
    .io_in_raddr(RAM_Block_18_io_in_raddr),
    .io_in_waddr(RAM_Block_18_io_in_waddr),
    .io_in_data_Re(RAM_Block_18_io_in_data_Re),
    .io_in_data_Im(RAM_Block_18_io_in_data_Im),
    .io_re(RAM_Block_18_io_re),
    .io_wr(RAM_Block_18_io_wr),
    .io_en(RAM_Block_18_io_en),
    .io_out_data_Re(RAM_Block_18_io_out_data_Re),
    .io_out_data_Im(RAM_Block_18_io_out_data_Im)
  );
  RAM_Block RAM_Block_19 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_19_clock),
    .io_in_raddr(RAM_Block_19_io_in_raddr),
    .io_in_waddr(RAM_Block_19_io_in_waddr),
    .io_in_data_Re(RAM_Block_19_io_in_data_Re),
    .io_in_data_Im(RAM_Block_19_io_in_data_Im),
    .io_re(RAM_Block_19_io_re),
    .io_wr(RAM_Block_19_io_wr),
    .io_en(RAM_Block_19_io_en),
    .io_out_data_Re(RAM_Block_19_io_out_data_Re),
    .io_out_data_Im(RAM_Block_19_io_out_data_Im)
  );
  RAM_Block RAM_Block_20 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_20_clock),
    .io_in_raddr(RAM_Block_20_io_in_raddr),
    .io_in_waddr(RAM_Block_20_io_in_waddr),
    .io_in_data_Re(RAM_Block_20_io_in_data_Re),
    .io_in_data_Im(RAM_Block_20_io_in_data_Im),
    .io_re(RAM_Block_20_io_re),
    .io_wr(RAM_Block_20_io_wr),
    .io_en(RAM_Block_20_io_en),
    .io_out_data_Re(RAM_Block_20_io_out_data_Re),
    .io_out_data_Im(RAM_Block_20_io_out_data_Im)
  );
  RAM_Block RAM_Block_21 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_21_clock),
    .io_in_raddr(RAM_Block_21_io_in_raddr),
    .io_in_waddr(RAM_Block_21_io_in_waddr),
    .io_in_data_Re(RAM_Block_21_io_in_data_Re),
    .io_in_data_Im(RAM_Block_21_io_in_data_Im),
    .io_re(RAM_Block_21_io_re),
    .io_wr(RAM_Block_21_io_wr),
    .io_en(RAM_Block_21_io_en),
    .io_out_data_Re(RAM_Block_21_io_out_data_Re),
    .io_out_data_Im(RAM_Block_21_io_out_data_Im)
  );
  RAM_Block RAM_Block_22 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_22_clock),
    .io_in_raddr(RAM_Block_22_io_in_raddr),
    .io_in_waddr(RAM_Block_22_io_in_waddr),
    .io_in_data_Re(RAM_Block_22_io_in_data_Re),
    .io_in_data_Im(RAM_Block_22_io_in_data_Im),
    .io_re(RAM_Block_22_io_re),
    .io_wr(RAM_Block_22_io_wr),
    .io_en(RAM_Block_22_io_en),
    .io_out_data_Re(RAM_Block_22_io_out_data_Re),
    .io_out_data_Im(RAM_Block_22_io_out_data_Im)
  );
  RAM_Block RAM_Block_23 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_23_clock),
    .io_in_raddr(RAM_Block_23_io_in_raddr),
    .io_in_waddr(RAM_Block_23_io_in_waddr),
    .io_in_data_Re(RAM_Block_23_io_in_data_Re),
    .io_in_data_Im(RAM_Block_23_io_in_data_Im),
    .io_re(RAM_Block_23_io_re),
    .io_wr(RAM_Block_23_io_wr),
    .io_en(RAM_Block_23_io_en),
    .io_out_data_Re(RAM_Block_23_io_out_data_Re),
    .io_out_data_Im(RAM_Block_23_io_out_data_Im)
  );
  RAM_Block RAM_Block_24 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_24_clock),
    .io_in_raddr(RAM_Block_24_io_in_raddr),
    .io_in_waddr(RAM_Block_24_io_in_waddr),
    .io_in_data_Re(RAM_Block_24_io_in_data_Re),
    .io_in_data_Im(RAM_Block_24_io_in_data_Im),
    .io_re(RAM_Block_24_io_re),
    .io_wr(RAM_Block_24_io_wr),
    .io_en(RAM_Block_24_io_en),
    .io_out_data_Re(RAM_Block_24_io_out_data_Re),
    .io_out_data_Im(RAM_Block_24_io_out_data_Im)
  );
  RAM_Block RAM_Block_25 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_25_clock),
    .io_in_raddr(RAM_Block_25_io_in_raddr),
    .io_in_waddr(RAM_Block_25_io_in_waddr),
    .io_in_data_Re(RAM_Block_25_io_in_data_Re),
    .io_in_data_Im(RAM_Block_25_io_in_data_Im),
    .io_re(RAM_Block_25_io_re),
    .io_wr(RAM_Block_25_io_wr),
    .io_en(RAM_Block_25_io_en),
    .io_out_data_Re(RAM_Block_25_io_out_data_Re),
    .io_out_data_Im(RAM_Block_25_io_out_data_Im)
  );
  RAM_Block RAM_Block_26 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_26_clock),
    .io_in_raddr(RAM_Block_26_io_in_raddr),
    .io_in_waddr(RAM_Block_26_io_in_waddr),
    .io_in_data_Re(RAM_Block_26_io_in_data_Re),
    .io_in_data_Im(RAM_Block_26_io_in_data_Im),
    .io_re(RAM_Block_26_io_re),
    .io_wr(RAM_Block_26_io_wr),
    .io_en(RAM_Block_26_io_en),
    .io_out_data_Re(RAM_Block_26_io_out_data_Re),
    .io_out_data_Im(RAM_Block_26_io_out_data_Im)
  );
  RAM_Block RAM_Block_27 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_27_clock),
    .io_in_raddr(RAM_Block_27_io_in_raddr),
    .io_in_waddr(RAM_Block_27_io_in_waddr),
    .io_in_data_Re(RAM_Block_27_io_in_data_Re),
    .io_in_data_Im(RAM_Block_27_io_in_data_Im),
    .io_re(RAM_Block_27_io_re),
    .io_wr(RAM_Block_27_io_wr),
    .io_en(RAM_Block_27_io_en),
    .io_out_data_Re(RAM_Block_27_io_out_data_Re),
    .io_out_data_Im(RAM_Block_27_io_out_data_Im)
  );
  RAM_Block RAM_Block_28 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_28_clock),
    .io_in_raddr(RAM_Block_28_io_in_raddr),
    .io_in_waddr(RAM_Block_28_io_in_waddr),
    .io_in_data_Re(RAM_Block_28_io_in_data_Re),
    .io_in_data_Im(RAM_Block_28_io_in_data_Im),
    .io_re(RAM_Block_28_io_re),
    .io_wr(RAM_Block_28_io_wr),
    .io_en(RAM_Block_28_io_en),
    .io_out_data_Re(RAM_Block_28_io_out_data_Re),
    .io_out_data_Im(RAM_Block_28_io_out_data_Im)
  );
  RAM_Block RAM_Block_29 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_29_clock),
    .io_in_raddr(RAM_Block_29_io_in_raddr),
    .io_in_waddr(RAM_Block_29_io_in_waddr),
    .io_in_data_Re(RAM_Block_29_io_in_data_Re),
    .io_in_data_Im(RAM_Block_29_io_in_data_Im),
    .io_re(RAM_Block_29_io_re),
    .io_wr(RAM_Block_29_io_wr),
    .io_en(RAM_Block_29_io_en),
    .io_out_data_Re(RAM_Block_29_io_out_data_Re),
    .io_out_data_Im(RAM_Block_29_io_out_data_Im)
  );
  RAM_Block RAM_Block_30 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_30_clock),
    .io_in_raddr(RAM_Block_30_io_in_raddr),
    .io_in_waddr(RAM_Block_30_io_in_waddr),
    .io_in_data_Re(RAM_Block_30_io_in_data_Re),
    .io_in_data_Im(RAM_Block_30_io_in_data_Im),
    .io_re(RAM_Block_30_io_re),
    .io_wr(RAM_Block_30_io_wr),
    .io_en(RAM_Block_30_io_en),
    .io_out_data_Re(RAM_Block_30_io_out_data_Re),
    .io_out_data_Im(RAM_Block_30_io_out_data_Im)
  );
  RAM_Block RAM_Block_31 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_31_clock),
    .io_in_raddr(RAM_Block_31_io_in_raddr),
    .io_in_waddr(RAM_Block_31_io_in_waddr),
    .io_in_data_Re(RAM_Block_31_io_in_data_Re),
    .io_in_data_Im(RAM_Block_31_io_in_data_Im),
    .io_re(RAM_Block_31_io_re),
    .io_wr(RAM_Block_31_io_wr),
    .io_en(RAM_Block_31_io_en),
    .io_out_data_Re(RAM_Block_31_io_out_data_Re),
    .io_out_data_Im(RAM_Block_31_io_out_data_Im)
  );
  PermutationModuleStreamed PermutationModuleStreamed ( // @[FFTDesigns.scala 2641:26]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_8_Re(PermutationModuleStreamed_io_in_8_Re),
    .io_in_8_Im(PermutationModuleStreamed_io_in_8_Im),
    .io_in_9_Re(PermutationModuleStreamed_io_in_9_Re),
    .io_in_9_Im(PermutationModuleStreamed_io_in_9_Im),
    .io_in_10_Re(PermutationModuleStreamed_io_in_10_Re),
    .io_in_10_Im(PermutationModuleStreamed_io_in_10_Im),
    .io_in_11_Re(PermutationModuleStreamed_io_in_11_Re),
    .io_in_11_Im(PermutationModuleStreamed_io_in_11_Im),
    .io_in_12_Re(PermutationModuleStreamed_io_in_12_Re),
    .io_in_12_Im(PermutationModuleStreamed_io_in_12_Im),
    .io_in_13_Re(PermutationModuleStreamed_io_in_13_Re),
    .io_in_13_Im(PermutationModuleStreamed_io_in_13_Im),
    .io_in_14_Re(PermutationModuleStreamed_io_in_14_Re),
    .io_in_14_Im(PermutationModuleStreamed_io_in_14_Im),
    .io_in_15_Re(PermutationModuleStreamed_io_in_15_Re),
    .io_in_15_Im(PermutationModuleStreamed_io_in_15_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_in_config_7(PermutationModuleStreamed_io_in_config_7),
    .io_in_config_8(PermutationModuleStreamed_io_in_config_8),
    .io_in_config_9(PermutationModuleStreamed_io_in_config_9),
    .io_in_config_10(PermutationModuleStreamed_io_in_config_10),
    .io_in_config_11(PermutationModuleStreamed_io_in_config_11),
    .io_in_config_12(PermutationModuleStreamed_io_in_config_12),
    .io_in_config_13(PermutationModuleStreamed_io_in_config_13),
    .io_in_config_14(PermutationModuleStreamed_io_in_config_14),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im),
    .io_out_8_Re(PermutationModuleStreamed_io_out_8_Re),
    .io_out_8_Im(PermutationModuleStreamed_io_out_8_Im),
    .io_out_9_Re(PermutationModuleStreamed_io_out_9_Re),
    .io_out_9_Im(PermutationModuleStreamed_io_out_9_Im),
    .io_out_10_Re(PermutationModuleStreamed_io_out_10_Re),
    .io_out_10_Im(PermutationModuleStreamed_io_out_10_Im),
    .io_out_11_Re(PermutationModuleStreamed_io_out_11_Re),
    .io_out_11_Im(PermutationModuleStreamed_io_out_11_Im),
    .io_out_12_Re(PermutationModuleStreamed_io_out_12_Re),
    .io_out_12_Im(PermutationModuleStreamed_io_out_12_Im),
    .io_out_13_Re(PermutationModuleStreamed_io_out_13_Re),
    .io_out_13_Im(PermutationModuleStreamed_io_out_13_Im),
    .io_out_14_Re(PermutationModuleStreamed_io_out_14_Re),
    .io_out_14_Im(PermutationModuleStreamed_io_out_14_Im),
    .io_out_15_Re(PermutationModuleStreamed_io_out_15_Re),
    .io_out_15_Im(PermutationModuleStreamed_io_out_15_Im)
  );
  M0_Config_ROM M0_Config_ROM ( // @[FFTDesigns.scala 2642:27]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7),
    .io_out_8(M0_Config_ROM_io_out_8),
    .io_out_9(M0_Config_ROM_io_out_9),
    .io_out_10(M0_Config_ROM_io_out_10),
    .io_out_11(M0_Config_ROM_io_out_11),
    .io_out_12(M0_Config_ROM_io_out_12),
    .io_out_13(M0_Config_ROM_io_out_13),
    .io_out_14(M0_Config_ROM_io_out_14),
    .io_out_15(M0_Config_ROM_io_out_15)
  );
  M1_Config_ROM M1_Config_ROM ( // @[FFTDesigns.scala 2643:27]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7),
    .io_out_8(M1_Config_ROM_io_out_8),
    .io_out_9(M1_Config_ROM_io_out_9),
    .io_out_10(M1_Config_ROM_io_out_10),
    .io_out_11(M1_Config_ROM_io_out_11),
    .io_out_12(M1_Config_ROM_io_out_12),
    .io_out_13(M1_Config_ROM_io_out_13),
    .io_out_14(M1_Config_ROM_io_out_14),
    .io_out_15(M1_Config_ROM_io_out_15)
  );
  Streaming_Permute_Config Streaming_Permute_Config ( // @[FFTDesigns.scala 2644:29]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6),
    .io_out_7(Streaming_Permute_Config_io_out_7),
    .io_out_8(Streaming_Permute_Config_io_out_8),
    .io_out_9(Streaming_Permute_Config_io_out_9),
    .io_out_10(Streaming_Permute_Config_io_out_10),
    .io_out_11(Streaming_Permute_Config_io_out_11),
    .io_out_12(Streaming_Permute_Config_io_out_12),
    .io_out_13(Streaming_Permute_Config_io_out_13),
    .io_out_14(Streaming_Permute_Config_io_out_14)
  );
  assign io_out_0_Re = RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_0_Im = RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Re = RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Im = RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Re = RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Im = RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Re = RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Im = RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Re = RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Im = RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Re = RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Im = RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Re = RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Im = RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Re = RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Im = RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_8_Re = RAM_Block_24_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_8_Im = RAM_Block_24_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_9_Re = RAM_Block_25_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_9_Im = RAM_Block_25_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_10_Re = RAM_Block_26_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_10_Im = RAM_Block_26_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_11_Re = RAM_Block_27_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_11_Im = RAM_Block_27_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_12_Re = RAM_Block_28_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_12_Im = RAM_Block_28_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_13_Re = RAM_Block_29_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_13_Im = RAM_Block_29_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_14_Re = RAM_Block_30_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_14_Im = RAM_Block_30_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_15_Re = RAM_Block_31_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_15_Im = RAM_Block_31_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = _GEN_6[1:0];
  assign RAM_Block_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_io_in_data_Re = io_in_0_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_in_data_Im = io_in_0_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = _GEN_19[1:0];
  assign RAM_Block_1_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_1_io_in_data_Re = io_in_1_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_in_data_Im = io_in_1_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = _GEN_32[1:0];
  assign RAM_Block_2_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_2_io_in_data_Re = io_in_2_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_in_data_Im = io_in_2_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = _GEN_45[1:0];
  assign RAM_Block_3_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_3_io_in_data_Re = io_in_3_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_in_data_Im = io_in_3_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = _GEN_58[1:0];
  assign RAM_Block_4_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_4_io_in_data_Re = io_in_4_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_in_data_Im = io_in_4_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = _GEN_71[1:0];
  assign RAM_Block_5_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_5_io_in_data_Re = io_in_5_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_in_data_Im = io_in_5_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = _GEN_84[1:0];
  assign RAM_Block_6_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_6_io_in_data_Re = io_in_6_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_in_data_Im = io_in_6_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = _GEN_97[1:0];
  assign RAM_Block_7_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_7_io_in_data_Re = io_in_7_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_in_data_Im = io_in_7_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = _GEN_110[1:0];
  assign RAM_Block_8_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_8_io_in_data_Re = io_in_8_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_8_io_in_data_Im = io_in_8_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = _GEN_123[1:0];
  assign RAM_Block_9_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_9_io_in_data_Re = io_in_9_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_9_io_in_data_Im = io_in_9_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = _GEN_136[1:0];
  assign RAM_Block_10_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_10_io_in_data_Re = io_in_10_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_10_io_in_data_Im = io_in_10_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = _GEN_149[1:0];
  assign RAM_Block_11_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_11_io_in_data_Re = io_in_11_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_11_io_in_data_Im = io_in_11_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = _GEN_162[1:0];
  assign RAM_Block_12_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_12_io_in_data_Re = io_in_12_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_12_io_in_data_Im = io_in_12_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = _GEN_175[1:0];
  assign RAM_Block_13_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_13_io_in_data_Re = io_in_13_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_13_io_in_data_Im = io_in_13_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = _GEN_188[1:0];
  assign RAM_Block_14_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_14_io_in_data_Re = io_in_14_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_14_io_in_data_Im = io_in_14_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = _GEN_201[1:0];
  assign RAM_Block_15_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_15_io_in_data_Re = io_in_15_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_15_io_in_data_Im = io_in_15_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_clock = clock;
  assign RAM_Block_16_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_16_io_in_waddr = _GEN_11[1:0];
  assign RAM_Block_16_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_16_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_16_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_clock = clock;
  assign RAM_Block_17_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_17_io_in_waddr = _GEN_24[1:0];
  assign RAM_Block_17_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_17_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_17_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_clock = clock;
  assign RAM_Block_18_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_18_io_in_waddr = _GEN_37[1:0];
  assign RAM_Block_18_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_18_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_18_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_clock = clock;
  assign RAM_Block_19_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_19_io_in_waddr = _GEN_50[1:0];
  assign RAM_Block_19_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_19_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_19_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_clock = clock;
  assign RAM_Block_20_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_20_io_in_waddr = _GEN_63[1:0];
  assign RAM_Block_20_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_20_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_20_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_clock = clock;
  assign RAM_Block_21_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_21_io_in_waddr = _GEN_76[1:0];
  assign RAM_Block_21_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_21_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_21_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_clock = clock;
  assign RAM_Block_22_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_22_io_in_waddr = _GEN_89[1:0];
  assign RAM_Block_22_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_22_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_22_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_clock = clock;
  assign RAM_Block_23_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_23_io_in_waddr = _GEN_102[1:0];
  assign RAM_Block_23_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_23_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_23_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_clock = clock;
  assign RAM_Block_24_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_24_io_in_waddr = _GEN_115[1:0];
  assign RAM_Block_24_io_in_data_Re = PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_24_io_in_data_Im = PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_24_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_clock = clock;
  assign RAM_Block_25_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_25_io_in_waddr = _GEN_128[1:0];
  assign RAM_Block_25_io_in_data_Re = PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_25_io_in_data_Im = PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_25_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_clock = clock;
  assign RAM_Block_26_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_26_io_in_waddr = _GEN_141[1:0];
  assign RAM_Block_26_io_in_data_Re = PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_26_io_in_data_Im = PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_26_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_clock = clock;
  assign RAM_Block_27_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_27_io_in_waddr = _GEN_154[1:0];
  assign RAM_Block_27_io_in_data_Re = PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_27_io_in_data_Im = PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_27_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_clock = clock;
  assign RAM_Block_28_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_28_io_in_waddr = _GEN_167[1:0];
  assign RAM_Block_28_io_in_data_Re = PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_28_io_in_data_Im = PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_28_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_clock = clock;
  assign RAM_Block_29_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_29_io_in_waddr = _GEN_180[1:0];
  assign RAM_Block_29_io_in_data_Re = PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_29_io_in_data_Im = PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_29_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_clock = clock;
  assign RAM_Block_30_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_30_io_in_waddr = _GEN_193[1:0];
  assign RAM_Block_30_io_in_data_Re = PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_30_io_in_data_Im = PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_30_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_clock = clock;
  assign RAM_Block_31_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_31_io_in_waddr = _GEN_206[1:0];
  assign RAM_Block_31_io_in_data_Re = PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_31_io_in_data_Im = PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_31_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_8_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_8_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_9_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_9_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_10_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_10_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_11_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_11_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_12_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_12_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_13_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_13_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_14_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_14_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_15_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_15_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_7 = Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_8 = Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_9 = Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_10 = Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_11 = Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_12 = Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_13 = Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_14 = Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign M0_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2694:22]
  assign M1_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2695:22]
  assign Streaming_Permute_Config_io_in_cnt = cnt; // @[FFTDesigns.scala 2696:24]
  always @(posedge clock) begin
    offset_switch <= _T_1 & _GEN_2; // @[FFTDesigns.scala 2646:30 2691:21]
    if (reset) begin // @[FFTDesigns.scala 2645:22]
      cnt <= 1'h0; // @[FFTDesigns.scala 2645:22]
    end else begin
      cnt <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module M1_Config_ROM_1(
  input        io_in_cnt,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2,
  output [1:0] io_out_3,
  output [1:0] io_out_4,
  output [1:0] io_out_5,
  output [1:0] io_out_6,
  output [1:0] io_out_7,
  output [1:0] io_out_8,
  output [1:0] io_out_9,
  output [1:0] io_out_10,
  output [1:0] io_out_11,
  output [1:0] io_out_12,
  output [1:0] io_out_13,
  output [1:0] io_out_14,
  output [1:0] io_out_15
);
  assign io_out_0 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_1 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_2 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_3 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_4 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_5 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_6 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_7 = io_in_cnt ? 2'h1 : 2'h0; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_8 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_9 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_10 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_11 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_12 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_13 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_14 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_15 = io_in_cnt ? 2'h0 : 2'h1; // @[FFTDesigns.scala 3250:{17,17}]
endmodule
module Streaming_Permute_Config_1(
  input        io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11,
  output [3:0] io_out_12,
  output [3:0] io_out_13,
  output [3:0] io_out_14
);
  assign io_out_0 = io_in_cnt ? 4'h8 : 4'h0; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_1 = io_in_cnt ? 4'h0 : 4'h8; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_2 = io_in_cnt ? 4'h9 : 4'h1; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_3 = io_in_cnt ? 4'h1 : 4'h9; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_4 = io_in_cnt ? 4'ha : 4'h2; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_5 = io_in_cnt ? 4'h2 : 4'ha; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_6 = io_in_cnt ? 4'hb : 4'h3; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_7 = io_in_cnt ? 4'h3 : 4'hb; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_8 = io_in_cnt ? 4'hc : 4'h4; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_9 = io_in_cnt ? 4'h4 : 4'hc; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_10 = io_in_cnt ? 4'hd : 4'h5; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_11 = io_in_cnt ? 4'h5 : 4'hd; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_12 = io_in_cnt ? 4'he : 4'h6; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_13 = io_in_cnt ? 4'h6 : 4'he; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_14 = io_in_cnt ? 4'hf : 4'h7; // @[FFTDesigns.scala 3273:{17,17}]
endmodule
module PermutationsWithStreaming_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [1:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_16_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_16_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_16_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_17_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_17_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_18_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_18_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_19_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_19_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_20_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_20_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_21_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_21_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_22_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_22_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_23_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_23_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_24_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_24_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_25_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_25_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_26_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_26_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_27_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_27_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_28_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_28_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_29_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_29_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_30_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_30_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_clock; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_31_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [1:0] RAM_Block_31_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_8_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_8_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_9_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_9_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_10_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_10_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_11_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_11_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_12_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_12_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_13_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_13_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_14_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_14_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_15_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_15_Im; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_7; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_8; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_9; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_10; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_11; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_12; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_13; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_14; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2641:26]
  wire  M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_8; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_9; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_10; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_11; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_12; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_13; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_14; // @[FFTDesigns.scala 2642:27]
  wire [1:0] M0_Config_ROM_io_out_15; // @[FFTDesigns.scala 2642:27]
  wire  M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_8; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_9; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_10; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_11; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_12; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_13; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_14; // @[FFTDesigns.scala 2643:27]
  wire [1:0] M1_Config_ROM_io_out_15; // @[FFTDesigns.scala 2643:27]
  wire  Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2644:29]
  reg  offset_switch; // @[FFTDesigns.scala 2627:28]
  wire [4:0] _T = {io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2628:19]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2628:26]
  reg  cnt; // @[FFTDesigns.scala 2645:22]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2649:26]
  wire  _GEN_1 = cnt ? 1'h0 : cnt + 1'h1; // @[FFTDesigns.scala 2647:32 2648:13 2651:13]
  wire  _GEN_2 = cnt ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2647:32 2649:23 2652:23]
  wire [2:0] _T_6 = 2'h2 * _offset_switch_T; // @[FFTDesigns.scala 2661:54]
  wire [2:0] _GEN_214 = {{1'd0}, M0_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_8 = _GEN_214 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_9 = 2'h2 * offset_switch; // @[FFTDesigns.scala 2662:41]
  wire [2:0] _GEN_215 = {{2'd0}, cnt}; // @[FFTDesigns.scala 2662:31]
  wire [2:0] _T_11 = _GEN_215 + _T_9; // @[FFTDesigns.scala 2662:31]
  wire [2:0] _T_15 = _GEN_215 + _T_6; // @[FFTDesigns.scala 2664:31]
  wire [2:0] _GEN_217 = {{1'd0}, M1_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_18 = _GEN_217 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_218 = {{1'd0}, M0_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_22 = _GEN_218 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_221 = {{1'd0}, M1_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_32 = _GEN_221 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_222 = {{1'd0}, M0_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_36 = _GEN_222 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_225 = {{1'd0}, M1_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_46 = _GEN_225 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_226 = {{1'd0}, M0_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_50 = _GEN_226 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_229 = {{1'd0}, M1_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_60 = _GEN_229 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_230 = {{1'd0}, M0_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_64 = _GEN_230 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_233 = {{1'd0}, M1_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_74 = _GEN_233 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_234 = {{1'd0}, M0_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_78 = _GEN_234 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_237 = {{1'd0}, M1_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_88 = _GEN_237 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_238 = {{1'd0}, M0_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_92 = _GEN_238 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_241 = {{1'd0}, M1_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_102 = _GEN_241 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_242 = {{1'd0}, M0_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_106 = _GEN_242 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_245 = {{1'd0}, M1_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_116 = _GEN_245 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_246 = {{1'd0}, M0_Config_ROM_io_out_8}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_120 = _GEN_246 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_249 = {{1'd0}, M1_Config_ROM_io_out_8}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_130 = _GEN_249 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_250 = {{1'd0}, M0_Config_ROM_io_out_9}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_134 = _GEN_250 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_253 = {{1'd0}, M1_Config_ROM_io_out_9}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_144 = _GEN_253 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_254 = {{1'd0}, M0_Config_ROM_io_out_10}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_148 = _GEN_254 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_257 = {{1'd0}, M1_Config_ROM_io_out_10}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_158 = _GEN_257 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_258 = {{1'd0}, M0_Config_ROM_io_out_11}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_162 = _GEN_258 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_261 = {{1'd0}, M1_Config_ROM_io_out_11}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_172 = _GEN_261 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_262 = {{1'd0}, M0_Config_ROM_io_out_12}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_176 = _GEN_262 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_265 = {{1'd0}, M1_Config_ROM_io_out_12}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_186 = _GEN_265 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_266 = {{1'd0}, M0_Config_ROM_io_out_13}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_190 = _GEN_266 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_269 = {{1'd0}, M1_Config_ROM_io_out_13}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_200 = _GEN_269 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_270 = {{1'd0}, M0_Config_ROM_io_out_14}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_204 = _GEN_270 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_273 = {{1'd0}, M1_Config_ROM_io_out_14}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_214 = _GEN_273 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _GEN_274 = {{1'd0}, M0_Config_ROM_io_out_15}; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _T_218 = _GEN_274 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [2:0] _GEN_277 = {{1'd0}, M1_Config_ROM_io_out_15}; // @[FFTDesigns.scala 2665:44]
  wire [2:0] _T_228 = _GEN_277 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire  _GEN_3 = _T_1 & _GEN_1; // @[FFTDesigns.scala 2646:30 2692:11]
  wire [2:0] _GEN_6 = _T_1 ? _T_8 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_7 = _T_1 ? _T_11 : 3'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  wire [2:0] _GEN_10 = _T_1 ? _T_15 : 3'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  wire [2:0] _GEN_11 = _T_1 ? _T_18 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_19 = _T_1 ? _T_22 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_24 = _T_1 ? _T_32 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_32 = _T_1 ? _T_36 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_37 = _T_1 ? _T_46 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_45 = _T_1 ? _T_50 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_50 = _T_1 ? _T_60 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_58 = _T_1 ? _T_64 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_63 = _T_1 ? _T_74 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_71 = _T_1 ? _T_78 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_76 = _T_1 ? _T_88 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_84 = _T_1 ? _T_92 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_89 = _T_1 ? _T_102 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_97 = _T_1 ? _T_106 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_102 = _T_1 ? _T_116 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_110 = _T_1 ? _T_120 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_115 = _T_1 ? _T_130 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_123 = _T_1 ? _T_134 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_128 = _T_1 ? _T_144 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_136 = _T_1 ? _T_148 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_141 = _T_1 ? _T_158 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_149 = _T_1 ? _T_162 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_154 = _T_1 ? _T_172 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_162 = _T_1 ? _T_176 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_167 = _T_1 ? _T_186 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_175 = _T_1 ? _T_190 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_180 = _T_1 ? _T_200 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_188 = _T_1 ? _T_204 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_193 = _T_1 ? _T_214 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  wire [2:0] _GEN_201 = _T_1 ? _T_218 : 3'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  wire [2:0] _GEN_206 = _T_1 ? _T_228 : 3'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  RAM_Block RAM_Block ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block RAM_Block_1 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block RAM_Block_2 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block RAM_Block_3 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block RAM_Block_4 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block RAM_Block_5 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block RAM_Block_6 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block RAM_Block_7 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block RAM_Block_8 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block RAM_Block_9 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block RAM_Block_10 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block RAM_Block_11 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block RAM_Block_12 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block RAM_Block_13 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block RAM_Block_14 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block RAM_Block_15 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  RAM_Block RAM_Block_16 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_16_clock),
    .io_in_raddr(RAM_Block_16_io_in_raddr),
    .io_in_waddr(RAM_Block_16_io_in_waddr),
    .io_in_data_Re(RAM_Block_16_io_in_data_Re),
    .io_in_data_Im(RAM_Block_16_io_in_data_Im),
    .io_re(RAM_Block_16_io_re),
    .io_wr(RAM_Block_16_io_wr),
    .io_en(RAM_Block_16_io_en),
    .io_out_data_Re(RAM_Block_16_io_out_data_Re),
    .io_out_data_Im(RAM_Block_16_io_out_data_Im)
  );
  RAM_Block RAM_Block_17 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_17_clock),
    .io_in_raddr(RAM_Block_17_io_in_raddr),
    .io_in_waddr(RAM_Block_17_io_in_waddr),
    .io_in_data_Re(RAM_Block_17_io_in_data_Re),
    .io_in_data_Im(RAM_Block_17_io_in_data_Im),
    .io_re(RAM_Block_17_io_re),
    .io_wr(RAM_Block_17_io_wr),
    .io_en(RAM_Block_17_io_en),
    .io_out_data_Re(RAM_Block_17_io_out_data_Re),
    .io_out_data_Im(RAM_Block_17_io_out_data_Im)
  );
  RAM_Block RAM_Block_18 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_18_clock),
    .io_in_raddr(RAM_Block_18_io_in_raddr),
    .io_in_waddr(RAM_Block_18_io_in_waddr),
    .io_in_data_Re(RAM_Block_18_io_in_data_Re),
    .io_in_data_Im(RAM_Block_18_io_in_data_Im),
    .io_re(RAM_Block_18_io_re),
    .io_wr(RAM_Block_18_io_wr),
    .io_en(RAM_Block_18_io_en),
    .io_out_data_Re(RAM_Block_18_io_out_data_Re),
    .io_out_data_Im(RAM_Block_18_io_out_data_Im)
  );
  RAM_Block RAM_Block_19 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_19_clock),
    .io_in_raddr(RAM_Block_19_io_in_raddr),
    .io_in_waddr(RAM_Block_19_io_in_waddr),
    .io_in_data_Re(RAM_Block_19_io_in_data_Re),
    .io_in_data_Im(RAM_Block_19_io_in_data_Im),
    .io_re(RAM_Block_19_io_re),
    .io_wr(RAM_Block_19_io_wr),
    .io_en(RAM_Block_19_io_en),
    .io_out_data_Re(RAM_Block_19_io_out_data_Re),
    .io_out_data_Im(RAM_Block_19_io_out_data_Im)
  );
  RAM_Block RAM_Block_20 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_20_clock),
    .io_in_raddr(RAM_Block_20_io_in_raddr),
    .io_in_waddr(RAM_Block_20_io_in_waddr),
    .io_in_data_Re(RAM_Block_20_io_in_data_Re),
    .io_in_data_Im(RAM_Block_20_io_in_data_Im),
    .io_re(RAM_Block_20_io_re),
    .io_wr(RAM_Block_20_io_wr),
    .io_en(RAM_Block_20_io_en),
    .io_out_data_Re(RAM_Block_20_io_out_data_Re),
    .io_out_data_Im(RAM_Block_20_io_out_data_Im)
  );
  RAM_Block RAM_Block_21 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_21_clock),
    .io_in_raddr(RAM_Block_21_io_in_raddr),
    .io_in_waddr(RAM_Block_21_io_in_waddr),
    .io_in_data_Re(RAM_Block_21_io_in_data_Re),
    .io_in_data_Im(RAM_Block_21_io_in_data_Im),
    .io_re(RAM_Block_21_io_re),
    .io_wr(RAM_Block_21_io_wr),
    .io_en(RAM_Block_21_io_en),
    .io_out_data_Re(RAM_Block_21_io_out_data_Re),
    .io_out_data_Im(RAM_Block_21_io_out_data_Im)
  );
  RAM_Block RAM_Block_22 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_22_clock),
    .io_in_raddr(RAM_Block_22_io_in_raddr),
    .io_in_waddr(RAM_Block_22_io_in_waddr),
    .io_in_data_Re(RAM_Block_22_io_in_data_Re),
    .io_in_data_Im(RAM_Block_22_io_in_data_Im),
    .io_re(RAM_Block_22_io_re),
    .io_wr(RAM_Block_22_io_wr),
    .io_en(RAM_Block_22_io_en),
    .io_out_data_Re(RAM_Block_22_io_out_data_Re),
    .io_out_data_Im(RAM_Block_22_io_out_data_Im)
  );
  RAM_Block RAM_Block_23 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_23_clock),
    .io_in_raddr(RAM_Block_23_io_in_raddr),
    .io_in_waddr(RAM_Block_23_io_in_waddr),
    .io_in_data_Re(RAM_Block_23_io_in_data_Re),
    .io_in_data_Im(RAM_Block_23_io_in_data_Im),
    .io_re(RAM_Block_23_io_re),
    .io_wr(RAM_Block_23_io_wr),
    .io_en(RAM_Block_23_io_en),
    .io_out_data_Re(RAM_Block_23_io_out_data_Re),
    .io_out_data_Im(RAM_Block_23_io_out_data_Im)
  );
  RAM_Block RAM_Block_24 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_24_clock),
    .io_in_raddr(RAM_Block_24_io_in_raddr),
    .io_in_waddr(RAM_Block_24_io_in_waddr),
    .io_in_data_Re(RAM_Block_24_io_in_data_Re),
    .io_in_data_Im(RAM_Block_24_io_in_data_Im),
    .io_re(RAM_Block_24_io_re),
    .io_wr(RAM_Block_24_io_wr),
    .io_en(RAM_Block_24_io_en),
    .io_out_data_Re(RAM_Block_24_io_out_data_Re),
    .io_out_data_Im(RAM_Block_24_io_out_data_Im)
  );
  RAM_Block RAM_Block_25 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_25_clock),
    .io_in_raddr(RAM_Block_25_io_in_raddr),
    .io_in_waddr(RAM_Block_25_io_in_waddr),
    .io_in_data_Re(RAM_Block_25_io_in_data_Re),
    .io_in_data_Im(RAM_Block_25_io_in_data_Im),
    .io_re(RAM_Block_25_io_re),
    .io_wr(RAM_Block_25_io_wr),
    .io_en(RAM_Block_25_io_en),
    .io_out_data_Re(RAM_Block_25_io_out_data_Re),
    .io_out_data_Im(RAM_Block_25_io_out_data_Im)
  );
  RAM_Block RAM_Block_26 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_26_clock),
    .io_in_raddr(RAM_Block_26_io_in_raddr),
    .io_in_waddr(RAM_Block_26_io_in_waddr),
    .io_in_data_Re(RAM_Block_26_io_in_data_Re),
    .io_in_data_Im(RAM_Block_26_io_in_data_Im),
    .io_re(RAM_Block_26_io_re),
    .io_wr(RAM_Block_26_io_wr),
    .io_en(RAM_Block_26_io_en),
    .io_out_data_Re(RAM_Block_26_io_out_data_Re),
    .io_out_data_Im(RAM_Block_26_io_out_data_Im)
  );
  RAM_Block RAM_Block_27 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_27_clock),
    .io_in_raddr(RAM_Block_27_io_in_raddr),
    .io_in_waddr(RAM_Block_27_io_in_waddr),
    .io_in_data_Re(RAM_Block_27_io_in_data_Re),
    .io_in_data_Im(RAM_Block_27_io_in_data_Im),
    .io_re(RAM_Block_27_io_re),
    .io_wr(RAM_Block_27_io_wr),
    .io_en(RAM_Block_27_io_en),
    .io_out_data_Re(RAM_Block_27_io_out_data_Re),
    .io_out_data_Im(RAM_Block_27_io_out_data_Im)
  );
  RAM_Block RAM_Block_28 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_28_clock),
    .io_in_raddr(RAM_Block_28_io_in_raddr),
    .io_in_waddr(RAM_Block_28_io_in_waddr),
    .io_in_data_Re(RAM_Block_28_io_in_data_Re),
    .io_in_data_Im(RAM_Block_28_io_in_data_Im),
    .io_re(RAM_Block_28_io_re),
    .io_wr(RAM_Block_28_io_wr),
    .io_en(RAM_Block_28_io_en),
    .io_out_data_Re(RAM_Block_28_io_out_data_Re),
    .io_out_data_Im(RAM_Block_28_io_out_data_Im)
  );
  RAM_Block RAM_Block_29 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_29_clock),
    .io_in_raddr(RAM_Block_29_io_in_raddr),
    .io_in_waddr(RAM_Block_29_io_in_waddr),
    .io_in_data_Re(RAM_Block_29_io_in_data_Re),
    .io_in_data_Im(RAM_Block_29_io_in_data_Im),
    .io_re(RAM_Block_29_io_re),
    .io_wr(RAM_Block_29_io_wr),
    .io_en(RAM_Block_29_io_en),
    .io_out_data_Re(RAM_Block_29_io_out_data_Re),
    .io_out_data_Im(RAM_Block_29_io_out_data_Im)
  );
  RAM_Block RAM_Block_30 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_30_clock),
    .io_in_raddr(RAM_Block_30_io_in_raddr),
    .io_in_waddr(RAM_Block_30_io_in_waddr),
    .io_in_data_Re(RAM_Block_30_io_in_data_Re),
    .io_in_data_Im(RAM_Block_30_io_in_data_Im),
    .io_re(RAM_Block_30_io_re),
    .io_wr(RAM_Block_30_io_wr),
    .io_en(RAM_Block_30_io_en),
    .io_out_data_Re(RAM_Block_30_io_out_data_Re),
    .io_out_data_Im(RAM_Block_30_io_out_data_Im)
  );
  RAM_Block RAM_Block_31 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_31_clock),
    .io_in_raddr(RAM_Block_31_io_in_raddr),
    .io_in_waddr(RAM_Block_31_io_in_waddr),
    .io_in_data_Re(RAM_Block_31_io_in_data_Re),
    .io_in_data_Im(RAM_Block_31_io_in_data_Im),
    .io_re(RAM_Block_31_io_re),
    .io_wr(RAM_Block_31_io_wr),
    .io_en(RAM_Block_31_io_en),
    .io_out_data_Re(RAM_Block_31_io_out_data_Re),
    .io_out_data_Im(RAM_Block_31_io_out_data_Im)
  );
  PermutationModuleStreamed PermutationModuleStreamed ( // @[FFTDesigns.scala 2641:26]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_8_Re(PermutationModuleStreamed_io_in_8_Re),
    .io_in_8_Im(PermutationModuleStreamed_io_in_8_Im),
    .io_in_9_Re(PermutationModuleStreamed_io_in_9_Re),
    .io_in_9_Im(PermutationModuleStreamed_io_in_9_Im),
    .io_in_10_Re(PermutationModuleStreamed_io_in_10_Re),
    .io_in_10_Im(PermutationModuleStreamed_io_in_10_Im),
    .io_in_11_Re(PermutationModuleStreamed_io_in_11_Re),
    .io_in_11_Im(PermutationModuleStreamed_io_in_11_Im),
    .io_in_12_Re(PermutationModuleStreamed_io_in_12_Re),
    .io_in_12_Im(PermutationModuleStreamed_io_in_12_Im),
    .io_in_13_Re(PermutationModuleStreamed_io_in_13_Re),
    .io_in_13_Im(PermutationModuleStreamed_io_in_13_Im),
    .io_in_14_Re(PermutationModuleStreamed_io_in_14_Re),
    .io_in_14_Im(PermutationModuleStreamed_io_in_14_Im),
    .io_in_15_Re(PermutationModuleStreamed_io_in_15_Re),
    .io_in_15_Im(PermutationModuleStreamed_io_in_15_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_in_config_7(PermutationModuleStreamed_io_in_config_7),
    .io_in_config_8(PermutationModuleStreamed_io_in_config_8),
    .io_in_config_9(PermutationModuleStreamed_io_in_config_9),
    .io_in_config_10(PermutationModuleStreamed_io_in_config_10),
    .io_in_config_11(PermutationModuleStreamed_io_in_config_11),
    .io_in_config_12(PermutationModuleStreamed_io_in_config_12),
    .io_in_config_13(PermutationModuleStreamed_io_in_config_13),
    .io_in_config_14(PermutationModuleStreamed_io_in_config_14),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im),
    .io_out_8_Re(PermutationModuleStreamed_io_out_8_Re),
    .io_out_8_Im(PermutationModuleStreamed_io_out_8_Im),
    .io_out_9_Re(PermutationModuleStreamed_io_out_9_Re),
    .io_out_9_Im(PermutationModuleStreamed_io_out_9_Im),
    .io_out_10_Re(PermutationModuleStreamed_io_out_10_Re),
    .io_out_10_Im(PermutationModuleStreamed_io_out_10_Im),
    .io_out_11_Re(PermutationModuleStreamed_io_out_11_Re),
    .io_out_11_Im(PermutationModuleStreamed_io_out_11_Im),
    .io_out_12_Re(PermutationModuleStreamed_io_out_12_Re),
    .io_out_12_Im(PermutationModuleStreamed_io_out_12_Im),
    .io_out_13_Re(PermutationModuleStreamed_io_out_13_Re),
    .io_out_13_Im(PermutationModuleStreamed_io_out_13_Im),
    .io_out_14_Re(PermutationModuleStreamed_io_out_14_Re),
    .io_out_14_Im(PermutationModuleStreamed_io_out_14_Im),
    .io_out_15_Re(PermutationModuleStreamed_io_out_15_Re),
    .io_out_15_Im(PermutationModuleStreamed_io_out_15_Im)
  );
  M0_Config_ROM M0_Config_ROM ( // @[FFTDesigns.scala 2642:27]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7),
    .io_out_8(M0_Config_ROM_io_out_8),
    .io_out_9(M0_Config_ROM_io_out_9),
    .io_out_10(M0_Config_ROM_io_out_10),
    .io_out_11(M0_Config_ROM_io_out_11),
    .io_out_12(M0_Config_ROM_io_out_12),
    .io_out_13(M0_Config_ROM_io_out_13),
    .io_out_14(M0_Config_ROM_io_out_14),
    .io_out_15(M0_Config_ROM_io_out_15)
  );
  M1_Config_ROM_1 M1_Config_ROM ( // @[FFTDesigns.scala 2643:27]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7),
    .io_out_8(M1_Config_ROM_io_out_8),
    .io_out_9(M1_Config_ROM_io_out_9),
    .io_out_10(M1_Config_ROM_io_out_10),
    .io_out_11(M1_Config_ROM_io_out_11),
    .io_out_12(M1_Config_ROM_io_out_12),
    .io_out_13(M1_Config_ROM_io_out_13),
    .io_out_14(M1_Config_ROM_io_out_14),
    .io_out_15(M1_Config_ROM_io_out_15)
  );
  Streaming_Permute_Config_1 Streaming_Permute_Config ( // @[FFTDesigns.scala 2644:29]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6),
    .io_out_7(Streaming_Permute_Config_io_out_7),
    .io_out_8(Streaming_Permute_Config_io_out_8),
    .io_out_9(Streaming_Permute_Config_io_out_9),
    .io_out_10(Streaming_Permute_Config_io_out_10),
    .io_out_11(Streaming_Permute_Config_io_out_11),
    .io_out_12(Streaming_Permute_Config_io_out_12),
    .io_out_13(Streaming_Permute_Config_io_out_13),
    .io_out_14(Streaming_Permute_Config_io_out_14)
  );
  assign io_out_0_Re = RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_0_Im = RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Re = RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Im = RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Re = RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Im = RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Re = RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Im = RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Re = RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Im = RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Re = RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Im = RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Re = RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Im = RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Re = RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Im = RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_8_Re = RAM_Block_24_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_8_Im = RAM_Block_24_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_9_Re = RAM_Block_25_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_9_Im = RAM_Block_25_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_10_Re = RAM_Block_26_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_10_Im = RAM_Block_26_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_11_Re = RAM_Block_27_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_11_Im = RAM_Block_27_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_12_Re = RAM_Block_28_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_12_Im = RAM_Block_28_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_13_Re = RAM_Block_29_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_13_Im = RAM_Block_29_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_14_Re = RAM_Block_30_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_14_Im = RAM_Block_30_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_15_Re = RAM_Block_31_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_15_Im = RAM_Block_31_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = _GEN_6[1:0];
  assign RAM_Block_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_io_in_data_Re = io_in_0_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_in_data_Im = io_in_0_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = _GEN_19[1:0];
  assign RAM_Block_1_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_1_io_in_data_Re = io_in_1_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_in_data_Im = io_in_1_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = _GEN_32[1:0];
  assign RAM_Block_2_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_2_io_in_data_Re = io_in_2_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_in_data_Im = io_in_2_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = _GEN_45[1:0];
  assign RAM_Block_3_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_3_io_in_data_Re = io_in_3_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_in_data_Im = io_in_3_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = _GEN_58[1:0];
  assign RAM_Block_4_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_4_io_in_data_Re = io_in_4_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_in_data_Im = io_in_4_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = _GEN_71[1:0];
  assign RAM_Block_5_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_5_io_in_data_Re = io_in_5_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_in_data_Im = io_in_5_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = _GEN_84[1:0];
  assign RAM_Block_6_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_6_io_in_data_Re = io_in_6_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_in_data_Im = io_in_6_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = _GEN_97[1:0];
  assign RAM_Block_7_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_7_io_in_data_Re = io_in_7_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_in_data_Im = io_in_7_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = _GEN_110[1:0];
  assign RAM_Block_8_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_8_io_in_data_Re = io_in_8_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_8_io_in_data_Im = io_in_8_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = _GEN_123[1:0];
  assign RAM_Block_9_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_9_io_in_data_Re = io_in_9_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_9_io_in_data_Im = io_in_9_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = _GEN_136[1:0];
  assign RAM_Block_10_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_10_io_in_data_Re = io_in_10_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_10_io_in_data_Im = io_in_10_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = _GEN_149[1:0];
  assign RAM_Block_11_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_11_io_in_data_Re = io_in_11_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_11_io_in_data_Im = io_in_11_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = _GEN_162[1:0];
  assign RAM_Block_12_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_12_io_in_data_Re = io_in_12_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_12_io_in_data_Im = io_in_12_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = _GEN_175[1:0];
  assign RAM_Block_13_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_13_io_in_data_Re = io_in_13_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_13_io_in_data_Im = io_in_13_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = _GEN_188[1:0];
  assign RAM_Block_14_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_14_io_in_data_Re = io_in_14_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_14_io_in_data_Im = io_in_14_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = _GEN_201[1:0];
  assign RAM_Block_15_io_in_waddr = _GEN_7[1:0];
  assign RAM_Block_15_io_in_data_Re = io_in_15_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_15_io_in_data_Im = io_in_15_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_clock = clock;
  assign RAM_Block_16_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_16_io_in_waddr = _GEN_11[1:0];
  assign RAM_Block_16_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_16_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_16_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_clock = clock;
  assign RAM_Block_17_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_17_io_in_waddr = _GEN_24[1:0];
  assign RAM_Block_17_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_17_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_17_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_clock = clock;
  assign RAM_Block_18_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_18_io_in_waddr = _GEN_37[1:0];
  assign RAM_Block_18_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_18_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_18_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_clock = clock;
  assign RAM_Block_19_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_19_io_in_waddr = _GEN_50[1:0];
  assign RAM_Block_19_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_19_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_19_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_clock = clock;
  assign RAM_Block_20_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_20_io_in_waddr = _GEN_63[1:0];
  assign RAM_Block_20_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_20_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_20_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_clock = clock;
  assign RAM_Block_21_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_21_io_in_waddr = _GEN_76[1:0];
  assign RAM_Block_21_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_21_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_21_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_clock = clock;
  assign RAM_Block_22_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_22_io_in_waddr = _GEN_89[1:0];
  assign RAM_Block_22_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_22_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_22_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_clock = clock;
  assign RAM_Block_23_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_23_io_in_waddr = _GEN_102[1:0];
  assign RAM_Block_23_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_23_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_23_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_clock = clock;
  assign RAM_Block_24_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_24_io_in_waddr = _GEN_115[1:0];
  assign RAM_Block_24_io_in_data_Re = PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_24_io_in_data_Im = PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_24_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_clock = clock;
  assign RAM_Block_25_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_25_io_in_waddr = _GEN_128[1:0];
  assign RAM_Block_25_io_in_data_Re = PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_25_io_in_data_Im = PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_25_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_clock = clock;
  assign RAM_Block_26_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_26_io_in_waddr = _GEN_141[1:0];
  assign RAM_Block_26_io_in_data_Re = PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_26_io_in_data_Im = PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_26_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_clock = clock;
  assign RAM_Block_27_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_27_io_in_waddr = _GEN_154[1:0];
  assign RAM_Block_27_io_in_data_Re = PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_27_io_in_data_Im = PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_27_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_clock = clock;
  assign RAM_Block_28_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_28_io_in_waddr = _GEN_167[1:0];
  assign RAM_Block_28_io_in_data_Re = PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_28_io_in_data_Im = PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_28_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_clock = clock;
  assign RAM_Block_29_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_29_io_in_waddr = _GEN_180[1:0];
  assign RAM_Block_29_io_in_data_Re = PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_29_io_in_data_Im = PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_29_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_clock = clock;
  assign RAM_Block_30_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_30_io_in_waddr = _GEN_193[1:0];
  assign RAM_Block_30_io_in_data_Re = PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_30_io_in_data_Im = PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_30_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_clock = clock;
  assign RAM_Block_31_io_in_raddr = _GEN_10[1:0];
  assign RAM_Block_31_io_in_waddr = _GEN_206[1:0];
  assign RAM_Block_31_io_in_data_Re = PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_31_io_in_data_Im = PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_31_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_8_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_8_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_9_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_9_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_10_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_10_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_11_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_11_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_12_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_12_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_13_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_13_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_14_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_14_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_15_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_15_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_7 = Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_8 = Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_9 = Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_10 = Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_11 = Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_12 = Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_13 = Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_14 = Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign M0_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2694:22]
  assign M1_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2695:22]
  assign Streaming_Permute_Config_io_in_cnt = cnt; // @[FFTDesigns.scala 2696:24]
  always @(posedge clock) begin
    offset_switch <= _T_1 & _GEN_2; // @[FFTDesigns.scala 2646:30 2691:21]
    if (reset) begin // @[FFTDesigns.scala 2645:22]
      cnt <= 1'h0; // @[FFTDesigns.scala 2645:22]
    end else begin
      cnt <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM(
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_9_Re,
  output [31:0] io_out_data_9_Im,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_11_Im,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_13_Im,
  output [31:0] io_out_data_15_Re,
  output [31:0] io_out_data_15_Im
);
  assign io_out_data_1_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_1_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_3_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_3_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_5_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_5_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_7_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_7_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_9_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_9_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_11_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_11_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_13_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_13_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_15_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_15_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
endmodule
module TwiddleFactorsStreamed(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] TwiddleFactorROM_io_in_addr; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_9_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_9_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_11_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_11_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_13_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_13_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_15_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_15_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] cmplx_adj_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_1_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_1_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_1_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_1_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_1_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_1_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_1_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_2_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_2_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_2_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_2_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_2_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_2_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_2_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_3_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_3_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_3_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_3_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_3_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_3_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_3_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_4_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_4_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_4_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_4_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_4_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_4_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_4_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_5_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_5_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_5_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_5_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_5_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_5_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_5_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_6_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_6_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_6_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_6_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_6_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_6_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_6_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_7_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_7_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_7_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_7_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_7_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_7_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_7_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_8_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_8_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_8_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_8_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_8_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_8_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_8_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_9_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_9_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_9_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_9_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_9_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_9_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_9_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_10_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_10_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_10_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_10_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_10_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_10_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_10_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_11_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_11_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_11_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_11_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_11_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_11_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_11_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_12_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_12_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_12_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_12_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_12_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_12_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_12_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_13_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_13_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_13_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_13_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_13_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_13_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_13_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_14_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_14_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_14_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_14_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_14_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_14_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_14_io_out_Im; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_15_io_in_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_15_io_in_Im; // @[FFTDesigns.scala 2146:30]
  wire [7:0] cmplx_adj_15_io_in_adj; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_15_io_is_neg; // @[FFTDesigns.scala 2146:30]
  wire  cmplx_adj_15_io_is_flip; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_15_io_out_Re; // @[FFTDesigns.scala 2146:30]
  wire [31:0] cmplx_adj_15_io_out_Im; // @[FFTDesigns.scala 2146:30]
  reg  cnt; // @[FFTDesigns.scala 2139:24]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2140:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2140:28]
  wire  _GEN_1 = cnt ? 1'h0 : cnt + 1'h1; // @[FFTDesigns.scala 2150:34 2151:15 2153:15]
  wire  _GEN_8 = TwiddleFactorROM_io_out_data_1_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_9 = TwiddleFactorROM_io_out_data_1_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_1_Re[31] :
    TwiddleFactorROM_io_out_data_1_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_16 = TwiddleFactorROM_io_out_data_3_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_17 = TwiddleFactorROM_io_out_data_3_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_3_Re[31] :
    TwiddleFactorROM_io_out_data_3_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_24 = TwiddleFactorROM_io_out_data_5_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_25 = TwiddleFactorROM_io_out_data_5_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_5_Re[31] :
    TwiddleFactorROM_io_out_data_5_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_32 = TwiddleFactorROM_io_out_data_7_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_33 = TwiddleFactorROM_io_out_data_7_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_7_Re[31] :
    TwiddleFactorROM_io_out_data_7_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_40 = TwiddleFactorROM_io_out_data_9_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_41 = TwiddleFactorROM_io_out_data_9_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_9_Re[31] :
    TwiddleFactorROM_io_out_data_9_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_48 = TwiddleFactorROM_io_out_data_11_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_49 = TwiddleFactorROM_io_out_data_11_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_11_Re[31] :
    TwiddleFactorROM_io_out_data_11_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_56 = TwiddleFactorROM_io_out_data_13_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_57 = TwiddleFactorROM_io_out_data_13_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_13_Re[31] :
    TwiddleFactorROM_io_out_data_13_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_64 = TwiddleFactorROM_io_out_data_15_Re[30:0] == 31'h3f800000 ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2158:92 2159:36 2166:36]
  wire  _GEN_65 = TwiddleFactorROM_io_out_data_15_Re[30:0] == 31'h3f800000 ? TwiddleFactorROM_io_out_data_15_Re[31] :
    TwiddleFactorROM_io_out_data_15_Im[31]; // @[FFTDesigns.scala 2158:92]
  wire  _GEN_66 = _T_1 & _GEN_1; // @[FFTDesigns.scala 2149:32 2175:13]
  reg [31:0] result_regs_0_0_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_0_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_1_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_1_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_2_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_2_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_3_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_3_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_4_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_4_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_5_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_5_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_6_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_6_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_7_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_7_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_8_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_8_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_9_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_9_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_10_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_10_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_11_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_11_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_12_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_12_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_13_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_13_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_14_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_14_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_15_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_0_15_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_0_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_0_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_1_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_1_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_2_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_2_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_3_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_3_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_4_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_4_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_5_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_5_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_6_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_6_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_7_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_7_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_8_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_8_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_9_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_9_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_10_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_10_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_11_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_11_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_12_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_12_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_13_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_13_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_14_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_14_Im; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_15_Re; // @[FFTDesigns.scala 2183:32]
  reg [31:0] result_regs_1_15_Im; // @[FFTDesigns.scala 2183:32]
  TwiddleFactorROM TwiddleFactorROM ( // @[FFTDesigns.scala 2098:26]
    .io_in_addr(TwiddleFactorROM_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_io_out_data_1_Im),
    .io_out_data_3_Re(TwiddleFactorROM_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_io_out_data_3_Im),
    .io_out_data_5_Re(TwiddleFactorROM_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_io_out_data_7_Im),
    .io_out_data_9_Re(TwiddleFactorROM_io_out_data_9_Re),
    .io_out_data_9_Im(TwiddleFactorROM_io_out_data_9_Im),
    .io_out_data_11_Re(TwiddleFactorROM_io_out_data_11_Re),
    .io_out_data_11_Im(TwiddleFactorROM_io_out_data_11_Im),
    .io_out_data_13_Re(TwiddleFactorROM_io_out_data_13_Re),
    .io_out_data_13_Im(TwiddleFactorROM_io_out_data_13_Im),
    .io_out_data_15_Re(TwiddleFactorROM_io_out_data_15_Re),
    .io_out_data_15_Im(TwiddleFactorROM_io_out_data_15_Im)
  );
  cmplx_adj cmplx_adj ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  cmplx_adj cmplx_adj_1 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_1_io_in_Re),
    .io_in_Im(cmplx_adj_1_io_in_Im),
    .io_in_adj(cmplx_adj_1_io_in_adj),
    .io_is_neg(cmplx_adj_1_io_is_neg),
    .io_is_flip(cmplx_adj_1_io_is_flip),
    .io_out_Re(cmplx_adj_1_io_out_Re),
    .io_out_Im(cmplx_adj_1_io_out_Im)
  );
  cmplx_adj cmplx_adj_2 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_2_io_in_Re),
    .io_in_Im(cmplx_adj_2_io_in_Im),
    .io_in_adj(cmplx_adj_2_io_in_adj),
    .io_is_neg(cmplx_adj_2_io_is_neg),
    .io_is_flip(cmplx_adj_2_io_is_flip),
    .io_out_Re(cmplx_adj_2_io_out_Re),
    .io_out_Im(cmplx_adj_2_io_out_Im)
  );
  cmplx_adj cmplx_adj_3 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_3_io_in_Re),
    .io_in_Im(cmplx_adj_3_io_in_Im),
    .io_in_adj(cmplx_adj_3_io_in_adj),
    .io_is_neg(cmplx_adj_3_io_is_neg),
    .io_is_flip(cmplx_adj_3_io_is_flip),
    .io_out_Re(cmplx_adj_3_io_out_Re),
    .io_out_Im(cmplx_adj_3_io_out_Im)
  );
  cmplx_adj cmplx_adj_4 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_4_io_in_Re),
    .io_in_Im(cmplx_adj_4_io_in_Im),
    .io_in_adj(cmplx_adj_4_io_in_adj),
    .io_is_neg(cmplx_adj_4_io_is_neg),
    .io_is_flip(cmplx_adj_4_io_is_flip),
    .io_out_Re(cmplx_adj_4_io_out_Re),
    .io_out_Im(cmplx_adj_4_io_out_Im)
  );
  cmplx_adj cmplx_adj_5 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_5_io_in_Re),
    .io_in_Im(cmplx_adj_5_io_in_Im),
    .io_in_adj(cmplx_adj_5_io_in_adj),
    .io_is_neg(cmplx_adj_5_io_is_neg),
    .io_is_flip(cmplx_adj_5_io_is_flip),
    .io_out_Re(cmplx_adj_5_io_out_Re),
    .io_out_Im(cmplx_adj_5_io_out_Im)
  );
  cmplx_adj cmplx_adj_6 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_6_io_in_Re),
    .io_in_Im(cmplx_adj_6_io_in_Im),
    .io_in_adj(cmplx_adj_6_io_in_adj),
    .io_is_neg(cmplx_adj_6_io_is_neg),
    .io_is_flip(cmplx_adj_6_io_is_flip),
    .io_out_Re(cmplx_adj_6_io_out_Re),
    .io_out_Im(cmplx_adj_6_io_out_Im)
  );
  cmplx_adj cmplx_adj_7 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_7_io_in_Re),
    .io_in_Im(cmplx_adj_7_io_in_Im),
    .io_in_adj(cmplx_adj_7_io_in_adj),
    .io_is_neg(cmplx_adj_7_io_is_neg),
    .io_is_flip(cmplx_adj_7_io_is_flip),
    .io_out_Re(cmplx_adj_7_io_out_Re),
    .io_out_Im(cmplx_adj_7_io_out_Im)
  );
  cmplx_adj cmplx_adj_8 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_8_io_in_Re),
    .io_in_Im(cmplx_adj_8_io_in_Im),
    .io_in_adj(cmplx_adj_8_io_in_adj),
    .io_is_neg(cmplx_adj_8_io_is_neg),
    .io_is_flip(cmplx_adj_8_io_is_flip),
    .io_out_Re(cmplx_adj_8_io_out_Re),
    .io_out_Im(cmplx_adj_8_io_out_Im)
  );
  cmplx_adj cmplx_adj_9 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_9_io_in_Re),
    .io_in_Im(cmplx_adj_9_io_in_Im),
    .io_in_adj(cmplx_adj_9_io_in_adj),
    .io_is_neg(cmplx_adj_9_io_is_neg),
    .io_is_flip(cmplx_adj_9_io_is_flip),
    .io_out_Re(cmplx_adj_9_io_out_Re),
    .io_out_Im(cmplx_adj_9_io_out_Im)
  );
  cmplx_adj cmplx_adj_10 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_10_io_in_Re),
    .io_in_Im(cmplx_adj_10_io_in_Im),
    .io_in_adj(cmplx_adj_10_io_in_adj),
    .io_is_neg(cmplx_adj_10_io_is_neg),
    .io_is_flip(cmplx_adj_10_io_is_flip),
    .io_out_Re(cmplx_adj_10_io_out_Re),
    .io_out_Im(cmplx_adj_10_io_out_Im)
  );
  cmplx_adj cmplx_adj_11 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_11_io_in_Re),
    .io_in_Im(cmplx_adj_11_io_in_Im),
    .io_in_adj(cmplx_adj_11_io_in_adj),
    .io_is_neg(cmplx_adj_11_io_is_neg),
    .io_is_flip(cmplx_adj_11_io_is_flip),
    .io_out_Re(cmplx_adj_11_io_out_Re),
    .io_out_Im(cmplx_adj_11_io_out_Im)
  );
  cmplx_adj cmplx_adj_12 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_12_io_in_Re),
    .io_in_Im(cmplx_adj_12_io_in_Im),
    .io_in_adj(cmplx_adj_12_io_in_adj),
    .io_is_neg(cmplx_adj_12_io_is_neg),
    .io_is_flip(cmplx_adj_12_io_is_flip),
    .io_out_Re(cmplx_adj_12_io_out_Re),
    .io_out_Im(cmplx_adj_12_io_out_Im)
  );
  cmplx_adj cmplx_adj_13 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_13_io_in_Re),
    .io_in_Im(cmplx_adj_13_io_in_Im),
    .io_in_adj(cmplx_adj_13_io_in_adj),
    .io_is_neg(cmplx_adj_13_io_is_neg),
    .io_is_flip(cmplx_adj_13_io_is_flip),
    .io_out_Re(cmplx_adj_13_io_out_Re),
    .io_out_Im(cmplx_adj_13_io_out_Im)
  );
  cmplx_adj cmplx_adj_14 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_14_io_in_Re),
    .io_in_Im(cmplx_adj_14_io_in_Im),
    .io_in_adj(cmplx_adj_14_io_in_adj),
    .io_is_neg(cmplx_adj_14_io_is_neg),
    .io_is_flip(cmplx_adj_14_io_is_flip),
    .io_out_Re(cmplx_adj_14_io_out_Re),
    .io_out_Im(cmplx_adj_14_io_out_Im)
  );
  cmplx_adj cmplx_adj_15 ( // @[FFTDesigns.scala 2146:30]
    .io_in_Re(cmplx_adj_15_io_in_Re),
    .io_in_Im(cmplx_adj_15_io_in_Im),
    .io_in_adj(cmplx_adj_15_io_in_adj),
    .io_is_neg(cmplx_adj_15_io_is_neg),
    .io_is_flip(cmplx_adj_15_io_is_flip),
    .io_out_Re(cmplx_adj_15_io_out_Re),
    .io_out_Im(cmplx_adj_15_io_out_Im)
  );
  assign io_out_0_Re = result_regs_1_0_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_0_Im = result_regs_1_0_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_1_Re = result_regs_1_1_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_1_Im = result_regs_1_1_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_2_Re = result_regs_1_2_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_2_Im = result_regs_1_2_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_3_Re = result_regs_1_3_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_3_Im = result_regs_1_3_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_4_Re = result_regs_1_4_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_4_Im = result_regs_1_4_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_5_Re = result_regs_1_5_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_5_Im = result_regs_1_5_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_6_Re = result_regs_1_6_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_6_Im = result_regs_1_6_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_7_Re = result_regs_1_7_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_7_Im = result_regs_1_7_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_8_Re = result_regs_1_8_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_8_Im = result_regs_1_8_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_9_Re = result_regs_1_9_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_9_Im = result_regs_1_9_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_10_Re = result_regs_1_10_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_10_Im = result_regs_1_10_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_11_Re = result_regs_1_11_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_11_Im = result_regs_1_11_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_12_Re = result_regs_1_12_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_12_Im = result_regs_1_12_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_13_Re = result_regs_1_13_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_13_Im = result_regs_1_13_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_14_Re = result_regs_1_14_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_14_Im = result_regs_1_14_Im; // @[FFTDesigns.scala 2193:14]
  assign io_out_15_Re = result_regs_1_15_Re; // @[FFTDesigns.scala 2193:14]
  assign io_out_15_Im = result_regs_1_15_Im; // @[FFTDesigns.scala 2193:14]
  assign TwiddleFactorROM_io_in_addr = {{4'd0}, cnt}; // @[FFTDesigns.scala 2194:24]
  assign cmplx_adj_io_in_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_io_in_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_io_in_adj = 8'h0;
  assign cmplx_adj_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_1_io_in_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_1_io_in_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_1_io_in_adj = 8'h0;
  assign cmplx_adj_1_io_is_neg = _T_1 & _GEN_9; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_1_io_is_flip = _T_1 & _GEN_8; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_2_io_in_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_2_io_in_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_2_io_in_adj = 8'h0;
  assign cmplx_adj_2_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_2_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_3_io_in_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_3_io_in_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_3_io_in_adj = 8'h0;
  assign cmplx_adj_3_io_is_neg = _T_1 & _GEN_17; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_3_io_is_flip = _T_1 & _GEN_16; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_4_io_in_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_4_io_in_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_4_io_in_adj = 8'h0;
  assign cmplx_adj_4_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_4_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_5_io_in_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_5_io_in_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_5_io_in_adj = 8'h0;
  assign cmplx_adj_5_io_is_neg = _T_1 & _GEN_25; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_5_io_is_flip = _T_1 & _GEN_24; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_6_io_in_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_6_io_in_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_6_io_in_adj = 8'h0;
  assign cmplx_adj_6_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_6_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_7_io_in_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_7_io_in_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_7_io_in_adj = 8'h0;
  assign cmplx_adj_7_io_is_neg = _T_1 & _GEN_33; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_7_io_is_flip = _T_1 & _GEN_32; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_8_io_in_Re = _T_1 ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_8_io_in_Im = _T_1 ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_8_io_in_adj = 8'h0;
  assign cmplx_adj_8_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_8_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_9_io_in_Re = _T_1 ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_9_io_in_Im = _T_1 ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_9_io_in_adj = 8'h0;
  assign cmplx_adj_9_io_is_neg = _T_1 & _GEN_41; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_9_io_is_flip = _T_1 & _GEN_40; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_10_io_in_Re = _T_1 ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_10_io_in_Im = _T_1 ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_10_io_in_adj = 8'h0;
  assign cmplx_adj_10_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_10_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_11_io_in_Re = _T_1 ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_11_io_in_Im = _T_1 ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_11_io_in_adj = 8'h0;
  assign cmplx_adj_11_io_is_neg = _T_1 & _GEN_49; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_11_io_is_flip = _T_1 & _GEN_48; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_12_io_in_Re = _T_1 ? io_in_12_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_12_io_in_Im = _T_1 ? io_in_12_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_12_io_in_adj = 8'h0;
  assign cmplx_adj_12_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_12_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_13_io_in_Re = _T_1 ? io_in_13_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_13_io_in_Im = _T_1 ? io_in_13_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_13_io_in_adj = 8'h0;
  assign cmplx_adj_13_io_is_neg = _T_1 & _GEN_57; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_13_io_is_flip = _T_1 & _GEN_56; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_14_io_in_Re = _T_1 ? io_in_14_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_14_io_in_Im = _T_1 ? io_in_14_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_14_io_in_adj = 8'h0;
  assign cmplx_adj_14_io_is_neg = 1'h0; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_14_io_is_flip = 1'h0; // @[FFTDesigns.scala 2149:32 2179:34]
  assign cmplx_adj_15_io_in_Re = _T_1 ? io_in_15_Re : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_15_io_in_Im = _T_1 ? io_in_15_Im : 32'h0; // @[FFTDesigns.scala 2149:32 2156:29 2177:29]
  assign cmplx_adj_15_io_in_adj = 8'h0;
  assign cmplx_adj_15_io_is_neg = _T_1 & _GEN_65; // @[FFTDesigns.scala 2149:32 2180:33]
  assign cmplx_adj_15_io_is_flip = _T_1 & _GEN_64; // @[FFTDesigns.scala 2149:32 2179:34]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2139:24]
      cnt <= 1'h0; // @[FFTDesigns.scala 2139:24]
    end else begin
      cnt <= _GEN_66;
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_0_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_0_Re <= cmplx_adj_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_0_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_0_Im <= cmplx_adj_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_1_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_1_Re <= cmplx_adj_1_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_1_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_1_Im <= cmplx_adj_1_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_2_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_2_Re <= cmplx_adj_2_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_2_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_2_Im <= cmplx_adj_2_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_3_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_3_Re <= cmplx_adj_3_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_3_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_3_Im <= cmplx_adj_3_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_4_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_4_Re <= cmplx_adj_4_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_4_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_4_Im <= cmplx_adj_4_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_5_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_5_Re <= cmplx_adj_5_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_5_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_5_Im <= cmplx_adj_5_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_6_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_6_Re <= cmplx_adj_6_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_6_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_6_Im <= cmplx_adj_6_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_7_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_7_Re <= cmplx_adj_7_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_7_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_7_Im <= cmplx_adj_7_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_8_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_8_Re <= cmplx_adj_8_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_8_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_8_Im <= cmplx_adj_8_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_9_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_9_Re <= cmplx_adj_9_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_9_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_9_Im <= cmplx_adj_9_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_10_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_10_Re <= cmplx_adj_10_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_10_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_10_Im <= cmplx_adj_10_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_11_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_11_Re <= cmplx_adj_11_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_11_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_11_Im <= cmplx_adj_11_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_12_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_12_Re <= cmplx_adj_12_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_12_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_12_Im <= cmplx_adj_12_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_13_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_13_Re <= cmplx_adj_13_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_13_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_13_Im <= cmplx_adj_13_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_14_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_14_Re <= cmplx_adj_14_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_14_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_14_Im <= cmplx_adj_14_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_15_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_15_Re <= cmplx_adj_15_io_out_Re; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_0_15_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_0_15_Im <= cmplx_adj_15_io_out_Im; // @[FFTDesigns.scala 2187:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_0_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_0_Re <= result_regs_0_0_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_0_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_0_Im <= result_regs_0_0_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_1_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_1_Re <= result_regs_0_1_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_1_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_1_Im <= result_regs_0_1_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_2_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_2_Re <= result_regs_0_2_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_2_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_2_Im <= result_regs_0_2_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_3_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_3_Re <= result_regs_0_3_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_3_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_3_Im <= result_regs_0_3_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_4_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_4_Re <= result_regs_0_4_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_4_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_4_Im <= result_regs_0_4_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_5_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_5_Re <= result_regs_0_5_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_5_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_5_Im <= result_regs_0_5_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_6_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_6_Re <= result_regs_0_6_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_6_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_6_Im <= result_regs_0_6_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_7_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_7_Re <= result_regs_0_7_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_7_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_7_Im <= result_regs_0_7_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_8_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_8_Re <= result_regs_0_8_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_8_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_8_Im <= result_regs_0_8_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_9_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_9_Re <= result_regs_0_9_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_9_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_9_Im <= result_regs_0_9_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_10_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_10_Re <= result_regs_0_10_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_10_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_10_Im <= result_regs_0_10_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_11_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_11_Re <= result_regs_0_11_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_11_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_11_Im <= result_regs_0_11_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_12_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_12_Re <= result_regs_0_12_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_12_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_12_Im <= result_regs_0_12_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_13_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_13_Re <= result_regs_0_13_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_13_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_13_Im <= result_regs_0_13_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_14_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_14_Re <= result_regs_0_14_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_14_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_14_Im <= result_regs_0_14_Im; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_15_Re <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_15_Re <= result_regs_0_15_Re; // @[FFTDesigns.scala 2190:26]
    end
    if (reset) begin // @[FFTDesigns.scala 2183:32]
      result_regs_1_15_Im <= 32'h0; // @[FFTDesigns.scala 2183:32]
    end else begin
      result_regs_1_15_Im <= result_regs_0_15_Im; // @[FFTDesigns.scala 2190:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  result_regs_0_0_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  result_regs_0_0_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  result_regs_0_1_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  result_regs_0_1_Im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  result_regs_0_2_Re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  result_regs_0_2_Im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  result_regs_0_3_Re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  result_regs_0_3_Im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  result_regs_0_4_Re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  result_regs_0_4_Im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  result_regs_0_5_Re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  result_regs_0_5_Im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  result_regs_0_6_Re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  result_regs_0_6_Im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  result_regs_0_7_Re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  result_regs_0_7_Im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  result_regs_0_8_Re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  result_regs_0_8_Im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  result_regs_0_9_Re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  result_regs_0_9_Im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  result_regs_0_10_Re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  result_regs_0_10_Im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  result_regs_0_11_Re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  result_regs_0_11_Im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  result_regs_0_12_Re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  result_regs_0_12_Im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  result_regs_0_13_Re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  result_regs_0_13_Im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  result_regs_0_14_Re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  result_regs_0_14_Im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  result_regs_0_15_Re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  result_regs_0_15_Im = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  result_regs_1_0_Re = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  result_regs_1_0_Im = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  result_regs_1_1_Re = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  result_regs_1_1_Im = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  result_regs_1_2_Re = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  result_regs_1_2_Im = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  result_regs_1_3_Re = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  result_regs_1_3_Im = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  result_regs_1_4_Re = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  result_regs_1_4_Im = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  result_regs_1_5_Re = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  result_regs_1_5_Im = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  result_regs_1_6_Re = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  result_regs_1_6_Im = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  result_regs_1_7_Re = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  result_regs_1_7_Im = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  result_regs_1_8_Re = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  result_regs_1_8_Im = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  result_regs_1_9_Re = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  result_regs_1_9_Im = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  result_regs_1_10_Re = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  result_regs_1_10_Im = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  result_regs_1_11_Re = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  result_regs_1_11_Im = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  result_regs_1_12_Re = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  result_regs_1_12_Im = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  result_regs_1_13_Re = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  result_regs_1_13_Im = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  result_regs_1_14_Re = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  result_regs_1_14_Im = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  result_regs_1_15_Re = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  result_regs_1_15_Im = _RAND_64[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_1(
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_9_Re,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_15_Re
);
  assign io_out_data_1_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_1_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_3_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_3_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_5_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_5_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_7_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_7_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_9_Re = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_11_Re = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_13_Re = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_15_Re = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[FFTDesigns.scala 2058:{25,25}]
endmodule
module FP_subber(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_clock; // @[FPArithmetic.scala 414:26]
  wire  FP_adder_reset; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_in_a; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_in_b; // @[FPArithmetic.scala 414:26]
  wire [31:0] FP_adder_io_out_s; // @[FPArithmetic.scala 414:26]
  wire  _adjusted_in_b_T_1 = ~io_in_b[31]; // @[FPArithmetic.scala 417:23]
  FP_adder FP_adder ( // @[FPArithmetic.scala 414:26]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  assign io_out_s = FP_adder_io_out_s; // @[FPArithmetic.scala 420:14]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = io_in_a; // @[FPArithmetic.scala 418:22]
  assign FP_adder_io_in_b = {_adjusted_in_b_T_1,io_in_b[30:0]}; // @[FPArithmetic.scala 417:39]
endmodule
module multiplier(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[Arithmetic.scala 84:23]
endmodule
module full_adder_162(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 58:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 58:34]
  wire [8:0] result = _result_T_1[8:0]; // @[Arithmetic.scala 57:22 58:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 59:23]
endmodule
module FP_multiplier(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] multiplier_io_in_a; // @[FPArithmetic.scala 488:28]
  wire [23:0] multiplier_io_in_b; // @[FPArithmetic.scala 488:28]
  wire [47:0] multiplier_io_out_s; // @[FPArithmetic.scala 488:28]
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 493:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 493:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 493:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 493:24]
  wire [7:0] complementN_io_in; // @[FPArithmetic.scala 499:29]
  wire [7:0] complementN_io_out; // @[FPArithmetic.scala 499:29]
  wire [7:0] adderN_io_in_a; // @[FPArithmetic.scala 503:24]
  wire [7:0] adderN_io_in_b; // @[FPArithmetic.scala 503:24]
  wire [7:0] adderN_io_out_s; // @[FPArithmetic.scala 503:24]
  wire  s_0 = io_in_a[31]; // @[FPArithmetic.scala 453:20]
  wire  s_1 = io_in_b[31]; // @[FPArithmetic.scala 454:20]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 458:62]
  wire [8:0] _GEN_13 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 458:34]
  wire [8:0] _GEN_0 = _GEN_13 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 458:68 459:14 461:14]
  wire [8:0] _GEN_14 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 463:34]
  wire [8:0] _GEN_1 = _GEN_14 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 463:68 464:14 466:14]
  wire [22:0] exp_check_0 = {{15'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 469:25 470:18]
  wire [22:0] _cond_holder_T_1 = exp_check_0 + 23'h1; // @[FPArithmetic.scala 474:34]
  wire [22:0] exp_check_1 = {{15'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 469:25 471:18]
  wire [22:0] _cond_holder_T_3 = 23'h7f - exp_check_1; // @[FPArithmetic.scala 474:80]
  wire [22:0] _cond_holder_T_4 = ~_cond_holder_T_3; // @[FPArithmetic.scala 474:42]
  wire [22:0] _cond_holder_T_6 = _cond_holder_T_1 + _cond_holder_T_4; // @[FPArithmetic.scala 474:40]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 478:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 479:23]
  wire  new_s = s_0 ^ s_1; // @[FPArithmetic.scala 510:19]
  wire [7:0] _new_exp_T_1 = adderN_io_out_s + 8'h1; // @[FPArithmetic.scala 521:34]
  wire [22:0] _cond_holder_T_8 = exp_check_0 + 23'h2; // @[FPArithmetic.scala 523:36]
  wire [22:0] _cond_holder_T_13 = _cond_holder_T_8 + _cond_holder_T_4; // @[FPArithmetic.scala 523:42]
  wire [23:0] _new_mant_T_2 = {multiplier_io_out_s[46:24], 1'h0}; // @[FPArithmetic.scala 529:73]
  wire [7:0] _GEN_2 = multiplier_io_out_s[47] ? _new_exp_T_1 : adderN_io_out_s; // @[FPArithmetic.scala 520:60 521:15 526:15]
  wire [22:0] cond_holder = multiplier_io_out_s[47] ? _cond_holder_T_13 : _cond_holder_T_6; // @[FPArithmetic.scala 520:60 523:19 528:19]
  wire [23:0] _GEN_5 = multiplier_io_out_s[47] ? {{1'd0}, multiplier_io_out_s[46:24]} : _new_mant_T_2; // @[FPArithmetic.scala 520:60 524:16 529:16]
  reg [31:0] reg_out_s; // @[FPArithmetic.scala 531:28]
  wire [22:0] _T_12 = ~cond_holder; // @[FPArithmetic.scala 533:51]
  wire [22:0] _T_14 = 23'h1 + _T_12; // @[FPArithmetic.scala 533:49]
  wire [22:0] _GEN_15 = {{14'd0}, _T_2}; // @[FPArithmetic.scala 533:42]
  wire [8:0] _GEN_6 = cond_holder > _GEN_15 ? _T_2 : {{1'd0}, _GEN_2}; // @[FPArithmetic.scala 538:61 539:15]
  wire [8:0] _GEN_9 = _GEN_15 >= _T_14 ? 9'h1 : _GEN_6; // @[FPArithmetic.scala 533:67 534:15]
  wire [7:0] new_exp = _GEN_9[7:0]; // @[FPArithmetic.scala 513:23]
  wire [23:0] _new_mant_T_4 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 540:45]
  wire [23:0] _GEN_7 = cond_holder > _GEN_15 ? _new_mant_T_4 : _GEN_5; // @[FPArithmetic.scala 538:61 540:16]
  wire [23:0] _GEN_10 = _GEN_15 >= _T_14 ? 24'h400000 : _GEN_7; // @[FPArithmetic.scala 533:67 535:16]
  wire [22:0] new_mant = _GEN_10[22:0]; // @[FPArithmetic.scala 515:24]
  wire [31:0] _reg_out_s_T_1 = {new_s,new_exp,new_mant}; // @[FPArithmetic.scala 536:37]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 457:19]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 457:19]
  multiplier multiplier ( // @[FPArithmetic.scala 488:28]
    .io_in_a(multiplier_io_in_a),
    .io_in_b(multiplier_io_in_b),
    .io_out_s(multiplier_io_out_s)
  );
  full_subber subber ( // @[FPArithmetic.scala 493:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complementN ( // @[FPArithmetic.scala 499:29]
    .io_in(complementN_io_in),
    .io_out(complementN_io_out)
  );
  full_adder_162 adderN ( // @[FPArithmetic.scala 503:24]
    .io_in_a(adderN_io_in_a),
    .io_in_b(adderN_io_in_b),
    .io_out_s(adderN_io_out_s)
  );
  assign io_out_s = reg_out_s; // @[FPArithmetic.scala 548:14]
  assign multiplier_io_in_a = {1'h1,frac_0}; // @[FPArithmetic.scala 483:24]
  assign multiplier_io_in_b = {1'h1,frac_1}; // @[FPArithmetic.scala 484:24]
  assign subber_io_in_a = 8'h7f; // @[FPArithmetic.scala 494:20]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 457:19]
  assign complementN_io_in = subber_io_out_s; // @[FPArithmetic.scala 500:23]
  assign adderN_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 457:19]
  assign adderN_io_in_b = complementN_io_out; // @[FPArithmetic.scala 505:20]
  always @(posedge clock) begin
    if (reset) begin // @[FPArithmetic.scala 531:28]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 531:28]
    end else if (exp_0 == 8'h0 | exp_1 == 8'h0) begin // @[FPArithmetic.scala 543:43]
      reg_out_s <= 32'h0; // @[FPArithmetic.scala 544:17]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FPArithmetic.scala 546:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_out_s = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMult(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_subber_clock; // @[FPComplex.scala 123:24]
  wire  FP_subber_reset; // @[FPComplex.scala 123:24]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 123:24]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 123:24]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 123:24]
  wire  FP_adder_clock; // @[FPComplex.scala 124:24]
  wire  FP_adder_reset; // @[FPComplex.scala 124:24]
  wire [31:0] FP_adder_io_in_a; // @[FPComplex.scala 124:24]
  wire [31:0] FP_adder_io_in_b; // @[FPComplex.scala 124:24]
  wire [31:0] FP_adder_io_out_s; // @[FPComplex.scala 124:24]
  wire  FP_multiplier_clock; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_reset; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_1_reset; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_2_clock; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_2_reset; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_2_io_in_a; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_2_io_in_b; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_2_io_out_s; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_3_clock; // @[FPComplex.scala 126:26]
  wire  FP_multiplier_3_reset; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_3_io_in_a; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_3_io_in_b; // @[FPComplex.scala 126:26]
  wire [31:0] FP_multiplier_3_io_out_s; // @[FPComplex.scala 126:26]
  FP_subber FP_subber ( // @[FPComplex.scala 123:24]
    .clock(FP_subber_clock),
    .reset(FP_subber_reset),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_adder FP_adder ( // @[FPComplex.scala 124:24]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 126:26]
    .clock(FP_multiplier_clock),
    .reset(FP_multiplier_reset),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 126:26]
    .clock(FP_multiplier_1_clock),
    .reset(FP_multiplier_1_reset),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  FP_multiplier FP_multiplier_2 ( // @[FPComplex.scala 126:26]
    .clock(FP_multiplier_2_clock),
    .reset(FP_multiplier_2_reset),
    .io_in_a(FP_multiplier_2_io_in_a),
    .io_in_b(FP_multiplier_2_io_in_b),
    .io_out_s(FP_multiplier_2_io_out_s)
  );
  FP_multiplier FP_multiplier_3 ( // @[FPComplex.scala 126:26]
    .clock(FP_multiplier_3_clock),
    .reset(FP_multiplier_3_reset),
    .io_in_a(FP_multiplier_3_io_in_a),
    .io_in_b(FP_multiplier_3_io_in_b),
    .io_out_s(FP_multiplier_3_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 141:17]
  assign io_out_s_Im = FP_adder_io_out_s; // @[FPComplex.scala 142:17]
  assign FP_subber_clock = clock;
  assign FP_subber_reset = reset;
  assign FP_subber_io_in_a = FP_multiplier_io_out_s; // @[FPComplex.scala 137:17]
  assign FP_subber_io_in_b = FP_multiplier_1_io_out_s; // @[FPComplex.scala 138:17]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = FP_multiplier_2_io_out_s; // @[FPComplex.scala 139:17]
  assign FP_adder_io_in_b = FP_multiplier_3_io_out_s; // @[FPComplex.scala 140:17]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_reset = reset;
  assign FP_multiplier_io_in_a = io_in_a_Re; // @[FPComplex.scala 129:28]
  assign FP_multiplier_io_in_b = io_in_b_Re; // @[FPComplex.scala 130:28]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_reset = reset;
  assign FP_multiplier_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 131:28]
  assign FP_multiplier_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 132:28]
  assign FP_multiplier_2_clock = clock;
  assign FP_multiplier_2_reset = reset;
  assign FP_multiplier_2_io_in_a = io_in_a_Re; // @[FPComplex.scala 133:28]
  assign FP_multiplier_2_io_in_b = io_in_b_Im; // @[FPComplex.scala 134:28]
  assign FP_multiplier_3_clock = clock;
  assign FP_multiplier_3_reset = reset;
  assign FP_multiplier_3_io_in_a = io_in_a_Im; // @[FPComplex.scala 135:28]
  assign FP_multiplier_3_io_in_b = io_in_b_Re; // @[FPComplex.scala 136:28]
endmodule
module TwiddleFactorsStreamed_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] TwiddleFactorROM_io_in_addr; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_9_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_11_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_13_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_15_Re; // @[FFTDesigns.scala 2098:26]
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_8_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_8_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_9_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_9_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_10_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_10_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_11_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_11_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_12_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_12_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_13_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_13_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_14_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_14_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_15_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_15_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  reg  cnt; // @[FFTDesigns.scala 2106:24]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2107:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2107:28]
  wire  _GEN_1 = cnt ? 1'h0 : cnt + 1'h1; // @[FFTDesigns.scala 2117:34 2118:15 2120:15]
  wire  _GEN_2 = _T_1 & _GEN_1; // @[FFTDesigns.scala 2116:32 2131:13]
  TwiddleFactorROM_1 TwiddleFactorROM ( // @[FFTDesigns.scala 2098:26]
    .io_in_addr(TwiddleFactorROM_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_io_out_data_1_Im),
    .io_out_data_3_Re(TwiddleFactorROM_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_io_out_data_3_Im),
    .io_out_data_5_Re(TwiddleFactorROM_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_io_out_data_7_Im),
    .io_out_data_9_Re(TwiddleFactorROM_io_out_data_9_Re),
    .io_out_data_11_Re(TwiddleFactorROM_io_out_data_11_Re),
    .io_out_data_13_Re(TwiddleFactorROM_io_out_data_13_Re),
    .io_out_data_15_Re(TwiddleFactorROM_io_out_data_15_Re)
  );
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_clock),
    .reset(FPComplexMult_reset),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_1_clock),
    .reset(FPComplexMult_1_reset),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_2_clock),
    .reset(FPComplexMult_2_reset),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_3_clock),
    .reset(FPComplexMult_3_reset),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_4_clock),
    .reset(FPComplexMult_4_reset),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_5_clock),
    .reset(FPComplexMult_5_reset),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_6_clock),
    .reset(FPComplexMult_6_reset),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_7_clock),
    .reset(FPComplexMult_7_reset),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_8 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_8_clock),
    .reset(FPComplexMult_8_reset),
    .io_in_a_Re(FPComplexMult_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_8_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_9 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_9_clock),
    .reset(FPComplexMult_9_reset),
    .io_in_a_Re(FPComplexMult_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_9_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_10 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_10_clock),
    .reset(FPComplexMult_10_reset),
    .io_in_a_Re(FPComplexMult_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_10_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_11 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_11_clock),
    .reset(FPComplexMult_11_reset),
    .io_in_a_Re(FPComplexMult_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_11_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_12 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_12_clock),
    .reset(FPComplexMult_12_reset),
    .io_in_a_Re(FPComplexMult_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_12_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_13 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_13_clock),
    .reset(FPComplexMult_13_reset),
    .io_in_a_Re(FPComplexMult_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_13_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_14 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_14_clock),
    .reset(FPComplexMult_14_reset),
    .io_in_a_Re(FPComplexMult_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_14_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_15 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_15_clock),
    .reset(FPComplexMult_15_reset),
    .io_in_a_Re(FPComplexMult_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_15_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_8_Re = FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_8_Im = FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_9_Re = FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_9_Im = FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_10_Re = FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_10_Im = FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_11_Re = FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_11_Im = FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_12_Re = FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_12_Im = FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_13_Re = FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_13_Im = FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_14_Re = FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_14_Im = FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_15_Re = FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_15_Im = FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign TwiddleFactorROM_io_in_addr = {{4'd0}, cnt}; // @[FFTDesigns.scala 2136:24]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_reset = reset;
  assign FPComplexMult_io_in_a_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_a_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_reset = reset;
  assign FPComplexMult_1_io_in_a_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_a_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_reset = reset;
  assign FPComplexMult_2_io_in_a_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_a_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_reset = reset;
  assign FPComplexMult_3_io_in_a_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_a_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_reset = reset;
  assign FPComplexMult_4_io_in_a_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_a_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_reset = reset;
  assign FPComplexMult_5_io_in_a_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_a_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_reset = reset;
  assign FPComplexMult_6_io_in_a_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_a_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_reset = reset;
  assign FPComplexMult_7_io_in_a_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_a_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_8_clock = clock;
  assign FPComplexMult_8_reset = reset;
  assign FPComplexMult_8_io_in_a_Re = _T_1 ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_8_io_in_a_Im = _T_1 ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_8_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_8_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_9_clock = clock;
  assign FPComplexMult_9_reset = reset;
  assign FPComplexMult_9_io_in_a_Re = _T_1 ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_9_io_in_a_Im = _T_1 ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_9_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_9_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_9_io_in_b_Im = _T_1 ? 32'hbf3504f2 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_10_clock = clock;
  assign FPComplexMult_10_reset = reset;
  assign FPComplexMult_10_io_in_a_Re = _T_1 ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_10_io_in_a_Im = _T_1 ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_10_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_10_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_11_clock = clock;
  assign FPComplexMult_11_reset = reset;
  assign FPComplexMult_11_io_in_a_Re = _T_1 ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_11_io_in_a_Im = _T_1 ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_11_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_11_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_11_io_in_b_Im = _T_1 ? 32'hbf3504f2 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_12_clock = clock;
  assign FPComplexMult_12_reset = reset;
  assign FPComplexMult_12_io_in_a_Re = _T_1 ? io_in_12_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_12_io_in_a_Im = _T_1 ? io_in_12_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_12_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_12_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_13_clock = clock;
  assign FPComplexMult_13_reset = reset;
  assign FPComplexMult_13_io_in_a_Re = _T_1 ? io_in_13_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_13_io_in_a_Im = _T_1 ? io_in_13_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_13_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_13_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_13_io_in_b_Im = _T_1 ? 32'hbf3504f2 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_14_clock = clock;
  assign FPComplexMult_14_reset = reset;
  assign FPComplexMult_14_io_in_a_Re = _T_1 ? io_in_14_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_14_io_in_a_Im = _T_1 ? io_in_14_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_14_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_14_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_15_clock = clock;
  assign FPComplexMult_15_reset = reset;
  assign FPComplexMult_15_io_in_a_Re = _T_1 ? io_in_15_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_15_io_in_a_Im = _T_1 ? io_in_15_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_15_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_15_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_15_io_in_b_Im = _T_1 ? 32'hbf3504f2 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2106:24]
      cnt <= 1'h0; // @[FFTDesigns.scala 2106:24]
    end else begin
      cnt <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_2(
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_9_Re,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_13_Im,
  output [31:0] io_out_data_15_Re,
  output [31:0] io_out_data_15_Im
);
  assign io_out_data_1_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_1_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_3_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_3_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_5_Re = io_in_addr[0] ? 32'hbec3ef14 : 32'h3f6c835e; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_5_Im = io_in_addr[0] ? 32'hbf6c835e : 32'hbec3ef14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_7_Re = io_in_addr[0] ? 32'hbec3ef14 : 32'h3f6c835e; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_7_Im = io_in_addr[0] ? 32'hbf6c835e : 32'hbec3ef14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_9_Re = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_11_Re = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_13_Re = io_in_addr[0] ? 32'hbf6c835e : 32'h3ec3ef14; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_13_Im = io_in_addr[0] ? 32'hbec3ef14 : 32'hbf6c835e; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_15_Re = io_in_addr[0] ? 32'hbf6c835e : 32'h3ec3ef14; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_15_Im = io_in_addr[0] ? 32'hbec3ef14 : 32'hbf6c835e; // @[FFTDesigns.scala 2059:{25,25}]
endmodule
module TwiddleFactorsStreamed_2(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] TwiddleFactorROM_io_in_addr; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_9_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_11_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_13_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_13_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_15_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_15_Im; // @[FFTDesigns.scala 2098:26]
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_8_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_8_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_9_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_9_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_10_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_10_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_11_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_11_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_12_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_12_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_13_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_13_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_14_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_14_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_15_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_15_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  reg  cnt; // @[FFTDesigns.scala 2106:24]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2107:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2107:28]
  wire  _GEN_1 = cnt ? 1'h0 : cnt + 1'h1; // @[FFTDesigns.scala 2117:34 2118:15 2120:15]
  wire  _GEN_2 = _T_1 & _GEN_1; // @[FFTDesigns.scala 2116:32 2131:13]
  TwiddleFactorROM_2 TwiddleFactorROM ( // @[FFTDesigns.scala 2098:26]
    .io_in_addr(TwiddleFactorROM_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_io_out_data_1_Im),
    .io_out_data_3_Re(TwiddleFactorROM_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_io_out_data_3_Im),
    .io_out_data_5_Re(TwiddleFactorROM_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_io_out_data_7_Im),
    .io_out_data_9_Re(TwiddleFactorROM_io_out_data_9_Re),
    .io_out_data_11_Re(TwiddleFactorROM_io_out_data_11_Re),
    .io_out_data_13_Re(TwiddleFactorROM_io_out_data_13_Re),
    .io_out_data_13_Im(TwiddleFactorROM_io_out_data_13_Im),
    .io_out_data_15_Re(TwiddleFactorROM_io_out_data_15_Re),
    .io_out_data_15_Im(TwiddleFactorROM_io_out_data_15_Im)
  );
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_clock),
    .reset(FPComplexMult_reset),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_1_clock),
    .reset(FPComplexMult_1_reset),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_2_clock),
    .reset(FPComplexMult_2_reset),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_3_clock),
    .reset(FPComplexMult_3_reset),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_4_clock),
    .reset(FPComplexMult_4_reset),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_5_clock),
    .reset(FPComplexMult_5_reset),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_6_clock),
    .reset(FPComplexMult_6_reset),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_7_clock),
    .reset(FPComplexMult_7_reset),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_8 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_8_clock),
    .reset(FPComplexMult_8_reset),
    .io_in_a_Re(FPComplexMult_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_8_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_9 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_9_clock),
    .reset(FPComplexMult_9_reset),
    .io_in_a_Re(FPComplexMult_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_9_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_10 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_10_clock),
    .reset(FPComplexMult_10_reset),
    .io_in_a_Re(FPComplexMult_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_10_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_11 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_11_clock),
    .reset(FPComplexMult_11_reset),
    .io_in_a_Re(FPComplexMult_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_11_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_12 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_12_clock),
    .reset(FPComplexMult_12_reset),
    .io_in_a_Re(FPComplexMult_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_12_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_13 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_13_clock),
    .reset(FPComplexMult_13_reset),
    .io_in_a_Re(FPComplexMult_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_13_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_14 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_14_clock),
    .reset(FPComplexMult_14_reset),
    .io_in_a_Re(FPComplexMult_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_14_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_15 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_15_clock),
    .reset(FPComplexMult_15_reset),
    .io_in_a_Re(FPComplexMult_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_15_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_8_Re = FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_8_Im = FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_9_Re = FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_9_Im = FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_10_Re = FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_10_Im = FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_11_Re = FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_11_Im = FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_12_Re = FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_12_Im = FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_13_Re = FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_13_Im = FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_14_Re = FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_14_Im = FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_15_Re = FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_15_Im = FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign TwiddleFactorROM_io_in_addr = {{4'd0}, cnt}; // @[FFTDesigns.scala 2136:24]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_reset = reset;
  assign FPComplexMult_io_in_a_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_a_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_reset = reset;
  assign FPComplexMult_1_io_in_a_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_a_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_reset = reset;
  assign FPComplexMult_2_io_in_a_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_a_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_reset = reset;
  assign FPComplexMult_3_io_in_a_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_a_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_reset = reset;
  assign FPComplexMult_4_io_in_a_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_a_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_reset = reset;
  assign FPComplexMult_5_io_in_a_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_a_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_reset = reset;
  assign FPComplexMult_6_io_in_a_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_a_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_reset = reset;
  assign FPComplexMult_7_io_in_a_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_a_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_8_clock = clock;
  assign FPComplexMult_8_reset = reset;
  assign FPComplexMult_8_io_in_a_Re = _T_1 ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_8_io_in_a_Im = _T_1 ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_8_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_8_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_9_clock = clock;
  assign FPComplexMult_9_reset = reset;
  assign FPComplexMult_9_io_in_a_Re = _T_1 ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_9_io_in_a_Im = _T_1 ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_9_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_9_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_9_io_in_b_Im = _T_1 ? 32'hbf3504f2 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_10_clock = clock;
  assign FPComplexMult_10_reset = reset;
  assign FPComplexMult_10_io_in_a_Re = _T_1 ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_10_io_in_a_Im = _T_1 ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_10_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_10_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_11_clock = clock;
  assign FPComplexMult_11_reset = reset;
  assign FPComplexMult_11_io_in_a_Re = _T_1 ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_11_io_in_a_Im = _T_1 ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_11_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_11_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_11_io_in_b_Im = _T_1 ? 32'hbf3504f2 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_12_clock = clock;
  assign FPComplexMult_12_reset = reset;
  assign FPComplexMult_12_io_in_a_Re = _T_1 ? io_in_12_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_12_io_in_a_Im = _T_1 ? io_in_12_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_12_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_12_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_13_clock = clock;
  assign FPComplexMult_13_reset = reset;
  assign FPComplexMult_13_io_in_a_Re = _T_1 ? io_in_13_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_13_io_in_a_Im = _T_1 ? io_in_13_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_13_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_13_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_13_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_13_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_14_clock = clock;
  assign FPComplexMult_14_reset = reset;
  assign FPComplexMult_14_io_in_a_Re = _T_1 ? io_in_14_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_14_io_in_a_Im = _T_1 ? io_in_14_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_14_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_14_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_15_clock = clock;
  assign FPComplexMult_15_reset = reset;
  assign FPComplexMult_15_io_in_a_Re = _T_1 ? io_in_15_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_15_io_in_a_Im = _T_1 ? io_in_15_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_15_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_15_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_15_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_15_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2106:24]
      cnt <= 1'h0; // @[FFTDesigns.scala 2106:24]
    end else begin
      cnt <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_3(
  input  [4:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_3_Re,
  output [31:0] io_out_data_3_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_9_Re,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_11_Im,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_13_Im,
  output [31:0] io_out_data_15_Re,
  output [31:0] io_out_data_15_Im
);
  assign io_out_data_1_Re = io_in_addr[0] ? 32'h248d3131 : 32'h3f800000; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_1_Im = io_in_addr[0] ? 32'hbf800000 : 32'h80800000; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_3_Re = io_in_addr[0] ? 32'hbe47c5c0 : 32'h3f7b14be; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_3_Im = io_in_addr[0] ? 32'hbf7b14be : 32'hbe47c5c0; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_5_Re = io_in_addr[0] ? 32'hbec3ef14 : 32'h3f6c835e; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_5_Im = io_in_addr[0] ? 32'hbf6c835e : 32'hbec3ef14; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_7_Re = io_in_addr[0] ? 32'hbf0e39d8 : 32'h3f54db30; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_7_Im = io_in_addr[0] ? 32'hbf54db30 : 32'hbf0e39d8; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_9_Re = io_in_addr[0] ? 32'hbf3504f2 : 32'h3f3504f2; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_11_Re = io_in_addr[0] ? 32'hbf54db30 : 32'h3f0e39d8; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_11_Im = io_in_addr[0] ? 32'hbf0e39d8 : 32'hbf54db30; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_13_Re = io_in_addr[0] ? 32'hbf6c835e : 32'h3ec3ef14; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_13_Im = io_in_addr[0] ? 32'hbec3ef14 : 32'hbf6c835e; // @[FFTDesigns.scala 2059:{25,25}]
  assign io_out_data_15_Re = io_in_addr[0] ? 32'hbf7b14be : 32'h3e47c5c0; // @[FFTDesigns.scala 2058:{25,25}]
  assign io_out_data_15_Im = io_in_addr[0] ? 32'hbe47c5c0 : 32'hbf7b14be; // @[FFTDesigns.scala 2059:{25,25}]
endmodule
module TwiddleFactorsStreamed_3(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] TwiddleFactorROM_io_in_addr; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_1_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_3_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_5_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_7_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_9_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_11_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_11_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_13_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_13_Im; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_15_Re; // @[FFTDesigns.scala 2098:26]
  wire [31:0] TwiddleFactorROM_io_out_data_15_Im; // @[FFTDesigns.scala 2098:26]
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_1_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_2_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_3_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_4_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_5_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_6_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_7_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_8_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_8_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_9_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_9_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_10_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_10_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_11_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_11_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_12_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_12_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_13_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_13_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_14_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_14_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_15_clock; // @[FFTDesigns.scala 2113:30]
  wire  FPComplexMult_15_reset; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_a_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_a_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_b_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_in_b_Im; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 2113:30]
  wire [31:0] FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 2113:30]
  reg  cnt; // @[FFTDesigns.scala 2106:24]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2107:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2107:28]
  wire  _GEN_1 = cnt ? 1'h0 : cnt + 1'h1; // @[FFTDesigns.scala 2117:34 2118:15 2120:15]
  wire  _GEN_2 = _T_1 & _GEN_1; // @[FFTDesigns.scala 2116:32 2131:13]
  TwiddleFactorROM_3 TwiddleFactorROM ( // @[FFTDesigns.scala 2098:26]
    .io_in_addr(TwiddleFactorROM_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_io_out_data_1_Im),
    .io_out_data_3_Re(TwiddleFactorROM_io_out_data_3_Re),
    .io_out_data_3_Im(TwiddleFactorROM_io_out_data_3_Im),
    .io_out_data_5_Re(TwiddleFactorROM_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_io_out_data_7_Im),
    .io_out_data_9_Re(TwiddleFactorROM_io_out_data_9_Re),
    .io_out_data_11_Re(TwiddleFactorROM_io_out_data_11_Re),
    .io_out_data_11_Im(TwiddleFactorROM_io_out_data_11_Im),
    .io_out_data_13_Re(TwiddleFactorROM_io_out_data_13_Re),
    .io_out_data_13_Im(TwiddleFactorROM_io_out_data_13_Im),
    .io_out_data_15_Re(TwiddleFactorROM_io_out_data_15_Re),
    .io_out_data_15_Im(TwiddleFactorROM_io_out_data_15_Im)
  );
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_clock),
    .reset(FPComplexMult_reset),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_1_clock),
    .reset(FPComplexMult_1_reset),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_2_clock),
    .reset(FPComplexMult_2_reset),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_3_clock),
    .reset(FPComplexMult_3_reset),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_4_clock),
    .reset(FPComplexMult_4_reset),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_5_clock),
    .reset(FPComplexMult_5_reset),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_6_clock),
    .reset(FPComplexMult_6_reset),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_7_clock),
    .reset(FPComplexMult_7_reset),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_8 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_8_clock),
    .reset(FPComplexMult_8_reset),
    .io_in_a_Re(FPComplexMult_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_8_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_9 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_9_clock),
    .reset(FPComplexMult_9_reset),
    .io_in_a_Re(FPComplexMult_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_9_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_10 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_10_clock),
    .reset(FPComplexMult_10_reset),
    .io_in_a_Re(FPComplexMult_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_10_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_11 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_11_clock),
    .reset(FPComplexMult_11_reset),
    .io_in_a_Re(FPComplexMult_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_11_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_12 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_12_clock),
    .reset(FPComplexMult_12_reset),
    .io_in_a_Re(FPComplexMult_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_12_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_13 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_13_clock),
    .reset(FPComplexMult_13_reset),
    .io_in_a_Re(FPComplexMult_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_13_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_14 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_14_clock),
    .reset(FPComplexMult_14_reset),
    .io_in_a_Re(FPComplexMult_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_14_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_15 ( // @[FFTDesigns.scala 2113:30]
    .clock(FPComplexMult_15_clock),
    .reset(FPComplexMult_15_reset),
    .io_in_a_Re(FPComplexMult_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_15_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_8_Re = FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_8_Im = FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_9_Re = FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_9_Im = FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_10_Re = FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_10_Im = FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_11_Re = FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_11_Im = FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_12_Re = FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_12_Im = FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_13_Re = FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_13_Im = FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_14_Re = FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_14_Im = FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign io_out_15_Re = FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 2134:19]
  assign io_out_15_Im = FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 2134:19]
  assign TwiddleFactorROM_io_in_addr = {{4'd0}, cnt}; // @[FFTDesigns.scala 2136:24]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_reset = reset;
  assign FPComplexMult_io_in_a_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_a_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_reset = reset;
  assign FPComplexMult_1_io_in_a_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_a_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_1_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_1_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_1_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_1_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_reset = reset;
  assign FPComplexMult_2_io_in_a_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_a_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_2_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_2_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_reset = reset;
  assign FPComplexMult_3_io_in_a_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_a_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_3_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_3_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_3_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_3_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_reset = reset;
  assign FPComplexMult_4_io_in_a_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_a_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_4_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_4_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_reset = reset;
  assign FPComplexMult_5_io_in_a_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_a_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_5_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_5_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_5_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_5_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_reset = reset;
  assign FPComplexMult_6_io_in_a_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_a_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_6_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_6_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_reset = reset;
  assign FPComplexMult_7_io_in_a_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_a_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_7_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_7_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_7_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_7_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_8_clock = clock;
  assign FPComplexMult_8_reset = reset;
  assign FPComplexMult_8_io_in_a_Re = _T_1 ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_8_io_in_a_Im = _T_1 ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_8_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_8_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_9_clock = clock;
  assign FPComplexMult_9_reset = reset;
  assign FPComplexMult_9_io_in_a_Re = _T_1 ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_9_io_in_a_Im = _T_1 ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_9_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_9_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_9_io_in_b_Im = _T_1 ? 32'hbf3504f2 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_10_clock = clock;
  assign FPComplexMult_10_reset = reset;
  assign FPComplexMult_10_io_in_a_Re = _T_1 ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_10_io_in_a_Im = _T_1 ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_10_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_10_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_11_clock = clock;
  assign FPComplexMult_11_reset = reset;
  assign FPComplexMult_11_io_in_a_Re = _T_1 ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_11_io_in_a_Im = _T_1 ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_11_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_11_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_11_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_11_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_12_clock = clock;
  assign FPComplexMult_12_reset = reset;
  assign FPComplexMult_12_io_in_a_Re = _T_1 ? io_in_12_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_12_io_in_a_Im = _T_1 ? io_in_12_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_12_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_12_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_13_clock = clock;
  assign FPComplexMult_13_reset = reset;
  assign FPComplexMult_13_io_in_a_Re = _T_1 ? io_in_13_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_13_io_in_a_Im = _T_1 ? io_in_13_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_13_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_13_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_13_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_13_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_14_clock = clock;
  assign FPComplexMult_14_reset = reset;
  assign FPComplexMult_14_io_in_a_Re = _T_1 ? io_in_14_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_14_io_in_a_Im = _T_1 ? io_in_14_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_14_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_14_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_15_clock = clock;
  assign FPComplexMult_15_reset = reset;
  assign FPComplexMult_15_io_in_a_Re = _T_1 ? io_in_15_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_15_io_in_a_Im = _T_1 ? io_in_15_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2123:31 2128:31]
  assign FPComplexMult_15_io_in_b_Re = _T_1 ? TwiddleFactorROM_io_out_data_15_Re : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  assign FPComplexMult_15_io_in_b_Im = _T_1 ? TwiddleFactorROM_io_out_data_15_Im : 32'h0; // @[FFTDesigns.scala 2116:32 2124:31 2129:31]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2106:24]
      cnt <= 1'h0; // @[FFTDesigns.scala 2106:24]
    end else begin
      cnt <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FFT_sr_v2_streaming_nrv(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_ready,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
`endif // RANDOMIZE_REG_INIT
  wire  DFT_r_v2_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_1_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_1_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_2_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_2_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_3_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_3_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_4_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_4_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_4_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_5_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_5_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_5_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_6_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_6_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_6_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_7_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_7_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_7_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_8_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_8_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_8_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_9_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_9_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_9_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_10_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_10_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_10_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_11_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_11_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_11_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_12_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_12_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_12_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_13_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_13_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_13_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_14_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_14_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_14_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_15_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_15_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_15_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_16_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_16_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_16_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_17_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_17_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_17_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_18_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_18_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_18_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_19_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_19_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_19_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_20_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_20_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_20_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_20_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_20_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_20_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_20_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_20_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_20_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_20_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_21_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_21_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_21_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_21_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_21_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_21_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_21_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_21_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_21_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_21_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_22_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_22_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_22_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_22_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_22_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_22_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_22_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_22_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_22_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_22_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_23_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_23_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_23_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_23_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_23_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_23_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_23_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_23_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_23_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_23_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_24_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_24_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_24_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_24_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_24_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_24_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_24_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_24_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_24_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_24_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_25_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_25_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_25_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_25_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_25_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_25_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_25_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_25_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_25_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_25_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_26_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_26_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_26_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_26_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_26_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_26_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_26_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_26_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_26_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_26_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_27_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_27_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_27_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_27_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_27_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_27_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_27_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_27_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_27_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_27_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_28_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_28_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_28_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_28_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_28_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_28_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_28_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_28_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_28_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_28_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_29_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_29_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_29_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_29_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_29_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_29_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_29_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_29_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_29_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_29_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_30_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_30_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_30_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_30_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_30_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_30_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_30_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_30_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_30_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_30_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_31_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_31_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_31_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_31_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_31_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_31_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_31_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_31_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_31_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_31_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_32_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_32_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_32_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_32_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_32_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_32_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_32_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_32_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_32_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_32_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_33_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_33_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_33_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_33_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_33_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_33_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_33_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_33_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_33_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_33_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_34_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_34_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_34_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_34_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_34_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_34_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_34_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_34_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_34_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_34_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_35_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_35_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_35_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_35_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_35_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_35_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_35_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_35_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_35_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_35_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_36_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_36_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_36_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_36_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_36_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_36_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_36_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_36_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_36_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_36_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_37_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_37_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_37_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_37_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_37_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_37_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_37_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_37_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_37_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_37_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_38_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_38_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_38_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_38_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_38_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_38_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_38_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_38_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_38_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_38_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_39_clock; // @[FFTDesigns.scala 5100:30]
  wire  DFT_r_v2_39_reset; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_39_io_in_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_39_io_in_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_39_io_in_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_39_io_in_1_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_39_io_out_0_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_39_io_out_0_Im; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_39_io_out_1_Re; // @[FFTDesigns.scala 5100:30]
  wire [31:0] DFT_r_v2_39_io_out_1_Im; // @[FFTDesigns.scala 5100:30]
  wire  PermutationsWithStreaming_clock; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_reset; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_0_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_0_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_1_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_1_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_2_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_2_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_3_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_3_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_4_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_4_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_5_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_5_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_6_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_6_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_7_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_7_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_8_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_8_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_9_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_9_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_10_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_10_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_11_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_11_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_12_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_12_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_13_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_13_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_14_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_14_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_15_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_in_15_Im; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_0; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_1; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_2; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_3; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_io_in_en_4; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_0_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_0_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_1_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_1_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_2_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_2_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_3_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_3_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_4_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_4_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_5_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_5_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_6_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_6_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_7_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_7_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_8_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_8_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_9_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_9_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_10_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_10_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_11_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_11_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_12_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_12_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_13_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_13_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_14_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_14_Im; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_15_Re; // @[FFTDesigns.scala 5107:30]
  wire [31:0] PermutationsWithStreaming_io_out_15_Im; // @[FFTDesigns.scala 5107:30]
  wire  PermutationsWithStreaming_1_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_in_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_1_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_1_io_out_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_in_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_2_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_2_io_out_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_in_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_3_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_3_io_out_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_in_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_4_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_4_io_out_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_clock; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_reset; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_in_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_0; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_1; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_2; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_3; // @[FFTDesigns.scala 5110:30]
  wire  PermutationsWithStreaming_5_io_in_en_4; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_0_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_0_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_1_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_1_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_2_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_2_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_3_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_3_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_4_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_4_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_5_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_5_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_6_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_6_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_7_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_7_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_8_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_8_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_9_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_9_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_10_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_10_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_11_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_11_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_12_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_12_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_13_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_13_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_14_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_14_Im; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_15_Re; // @[FFTDesigns.scala 5110:30]
  wire [31:0] PermutationsWithStreaming_5_io_out_15_Im; // @[FFTDesigns.scala 5110:30]
  wire  TwiddleFactorsStreamed_clock; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_reset; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_7_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_8_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_8_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_9_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_9_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_10_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_10_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_11_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_11_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_12_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_12_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_13_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_13_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_14_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_14_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_15_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_in_15_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_io_in_en_0; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_io_in_en_1; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_7_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_8_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_8_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_9_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_9_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_10_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_10_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_11_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_11_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_12_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_12_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_13_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_13_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_14_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_14_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_15_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_io_out_15_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_1_clock; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_1_reset; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_7_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_8_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_8_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_9_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_9_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_10_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_10_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_11_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_11_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_12_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_12_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_13_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_13_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_14_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_14_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_15_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_in_15_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_1_io_in_en_0; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_1_io_in_en_1; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_7_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_8_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_8_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_9_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_9_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_10_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_10_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_11_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_11_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_12_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_12_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_13_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_13_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_14_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_14_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_15_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_1_io_out_15_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_2_clock; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_2_reset; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_7_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_8_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_8_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_9_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_9_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_10_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_10_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_11_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_11_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_12_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_12_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_13_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_13_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_14_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_14_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_15_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_in_15_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_2_io_in_en_0; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_2_io_in_en_1; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_7_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_8_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_8_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_9_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_9_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_10_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_10_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_11_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_11_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_12_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_12_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_13_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_13_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_14_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_14_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_15_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_2_io_out_15_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_3_clock; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_3_reset; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_7_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_8_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_8_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_9_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_9_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_10_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_10_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_11_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_11_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_12_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_12_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_13_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_13_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_14_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_14_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_15_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_in_15_Im; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_3_io_in_en_0; // @[FFTDesigns.scala 5115:28]
  wire  TwiddleFactorsStreamed_3_io_in_en_1; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_0_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_0_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_1_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_1_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_2_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_2_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_3_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_3_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_4_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_4_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_5_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_5_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_6_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_6_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_7_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_7_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_8_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_8_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_9_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_9_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_10_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_10_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_11_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_11_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_12_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_12_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_13_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_13_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_14_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_14_Im; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_15_Re; // @[FFTDesigns.scala 5115:28]
  wire [31:0] TwiddleFactorsStreamed_3_io_out_15_Im; // @[FFTDesigns.scala 5115:28]
  reg  DFT_regdelays_0_0; // @[FFTDesigns.scala 5094:32]
  reg  DFT_regdelays_1_0; // @[FFTDesigns.scala 5094:32]
  reg  DFT_regdelays_2_0; // @[FFTDesigns.scala 5094:32]
  reg  DFT_regdelays_3_0; // @[FFTDesigns.scala 5094:32]
  reg  DFT_regdelays_4_0; // @[FFTDesigns.scala 5094:32]
  reg  Twid_regdelays_0_0; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_0_1; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_1_0; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_1_1; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_2_0; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_2_1; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_3_0; // @[FFTDesigns.scala 5095:33]
  reg  Twid_regdelays_3_1; // @[FFTDesigns.scala 5095:33]
  reg  Perm_regdelays_0_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_0_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_1_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_2_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_3_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_4_3; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_0; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_1; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_2; // @[FFTDesigns.scala 5096:33]
  reg  Perm_regdelays_5_3; // @[FFTDesigns.scala 5096:33]
  DFT_r_v2 DFT_r_v2 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_clock),
    .reset(DFT_r_v2_reset),
    .io_in_0_Re(DFT_r_v2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_1 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_1_clock),
    .reset(DFT_r_v2_1_reset),
    .io_in_0_Re(DFT_r_v2_1_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_1_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_1_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_1_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_1_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_1_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_1_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_1_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_2 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_2_clock),
    .reset(DFT_r_v2_2_reset),
    .io_in_0_Re(DFT_r_v2_2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_2_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_2_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_3 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_3_clock),
    .reset(DFT_r_v2_3_reset),
    .io_in_0_Re(DFT_r_v2_3_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_3_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_3_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_3_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_3_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_3_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_3_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_3_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_4 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_4_clock),
    .reset(DFT_r_v2_4_reset),
    .io_in_0_Re(DFT_r_v2_4_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_4_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_4_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_4_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_4_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_4_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_4_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_4_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_5 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_5_clock),
    .reset(DFT_r_v2_5_reset),
    .io_in_0_Re(DFT_r_v2_5_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_5_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_5_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_5_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_5_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_5_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_5_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_5_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_6 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_6_clock),
    .reset(DFT_r_v2_6_reset),
    .io_in_0_Re(DFT_r_v2_6_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_6_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_6_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_6_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_6_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_6_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_6_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_6_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_7 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_7_clock),
    .reset(DFT_r_v2_7_reset),
    .io_in_0_Re(DFT_r_v2_7_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_7_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_7_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_7_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_7_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_7_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_7_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_7_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_8 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_8_clock),
    .reset(DFT_r_v2_8_reset),
    .io_in_0_Re(DFT_r_v2_8_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_8_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_8_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_8_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_8_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_8_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_8_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_8_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_9 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_9_clock),
    .reset(DFT_r_v2_9_reset),
    .io_in_0_Re(DFT_r_v2_9_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_9_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_9_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_9_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_9_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_9_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_9_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_9_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_10 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_10_clock),
    .reset(DFT_r_v2_10_reset),
    .io_in_0_Re(DFT_r_v2_10_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_10_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_10_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_10_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_10_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_10_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_10_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_10_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_11 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_11_clock),
    .reset(DFT_r_v2_11_reset),
    .io_in_0_Re(DFT_r_v2_11_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_11_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_11_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_11_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_11_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_11_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_11_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_11_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_12 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_12_clock),
    .reset(DFT_r_v2_12_reset),
    .io_in_0_Re(DFT_r_v2_12_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_12_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_12_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_12_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_12_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_12_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_12_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_12_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_13 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_13_clock),
    .reset(DFT_r_v2_13_reset),
    .io_in_0_Re(DFT_r_v2_13_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_13_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_13_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_13_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_13_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_13_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_13_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_13_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_14 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_14_clock),
    .reset(DFT_r_v2_14_reset),
    .io_in_0_Re(DFT_r_v2_14_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_14_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_14_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_14_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_14_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_14_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_14_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_14_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_15 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_15_clock),
    .reset(DFT_r_v2_15_reset),
    .io_in_0_Re(DFT_r_v2_15_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_15_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_15_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_15_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_15_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_15_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_15_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_15_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_16 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_16_clock),
    .reset(DFT_r_v2_16_reset),
    .io_in_0_Re(DFT_r_v2_16_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_16_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_16_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_16_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_16_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_16_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_16_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_16_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_17 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_17_clock),
    .reset(DFT_r_v2_17_reset),
    .io_in_0_Re(DFT_r_v2_17_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_17_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_17_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_17_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_17_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_17_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_17_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_17_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_18 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_18_clock),
    .reset(DFT_r_v2_18_reset),
    .io_in_0_Re(DFT_r_v2_18_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_18_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_18_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_18_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_18_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_18_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_18_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_18_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_19 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_19_clock),
    .reset(DFT_r_v2_19_reset),
    .io_in_0_Re(DFT_r_v2_19_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_19_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_19_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_19_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_19_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_19_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_19_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_19_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_20 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_20_clock),
    .reset(DFT_r_v2_20_reset),
    .io_in_0_Re(DFT_r_v2_20_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_20_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_20_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_20_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_20_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_20_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_20_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_20_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_21 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_21_clock),
    .reset(DFT_r_v2_21_reset),
    .io_in_0_Re(DFT_r_v2_21_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_21_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_21_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_21_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_21_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_21_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_21_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_21_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_22 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_22_clock),
    .reset(DFT_r_v2_22_reset),
    .io_in_0_Re(DFT_r_v2_22_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_22_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_22_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_22_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_22_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_22_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_22_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_22_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_23 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_23_clock),
    .reset(DFT_r_v2_23_reset),
    .io_in_0_Re(DFT_r_v2_23_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_23_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_23_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_23_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_23_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_23_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_23_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_23_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_24 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_24_clock),
    .reset(DFT_r_v2_24_reset),
    .io_in_0_Re(DFT_r_v2_24_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_24_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_24_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_24_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_24_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_24_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_24_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_24_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_25 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_25_clock),
    .reset(DFT_r_v2_25_reset),
    .io_in_0_Re(DFT_r_v2_25_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_25_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_25_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_25_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_25_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_25_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_25_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_25_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_26 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_26_clock),
    .reset(DFT_r_v2_26_reset),
    .io_in_0_Re(DFT_r_v2_26_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_26_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_26_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_26_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_26_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_26_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_26_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_26_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_27 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_27_clock),
    .reset(DFT_r_v2_27_reset),
    .io_in_0_Re(DFT_r_v2_27_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_27_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_27_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_27_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_27_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_27_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_27_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_27_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_28 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_28_clock),
    .reset(DFT_r_v2_28_reset),
    .io_in_0_Re(DFT_r_v2_28_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_28_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_28_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_28_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_28_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_28_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_28_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_28_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_29 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_29_clock),
    .reset(DFT_r_v2_29_reset),
    .io_in_0_Re(DFT_r_v2_29_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_29_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_29_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_29_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_29_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_29_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_29_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_29_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_30 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_30_clock),
    .reset(DFT_r_v2_30_reset),
    .io_in_0_Re(DFT_r_v2_30_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_30_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_30_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_30_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_30_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_30_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_30_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_30_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_31 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_31_clock),
    .reset(DFT_r_v2_31_reset),
    .io_in_0_Re(DFT_r_v2_31_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_31_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_31_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_31_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_31_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_31_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_31_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_31_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_32 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_32_clock),
    .reset(DFT_r_v2_32_reset),
    .io_in_0_Re(DFT_r_v2_32_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_32_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_32_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_32_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_32_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_32_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_32_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_32_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_33 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_33_clock),
    .reset(DFT_r_v2_33_reset),
    .io_in_0_Re(DFT_r_v2_33_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_33_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_33_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_33_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_33_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_33_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_33_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_33_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_34 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_34_clock),
    .reset(DFT_r_v2_34_reset),
    .io_in_0_Re(DFT_r_v2_34_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_34_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_34_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_34_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_34_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_34_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_34_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_34_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_35 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_35_clock),
    .reset(DFT_r_v2_35_reset),
    .io_in_0_Re(DFT_r_v2_35_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_35_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_35_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_35_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_35_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_35_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_35_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_35_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_36 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_36_clock),
    .reset(DFT_r_v2_36_reset),
    .io_in_0_Re(DFT_r_v2_36_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_36_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_36_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_36_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_36_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_36_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_36_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_36_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_37 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_37_clock),
    .reset(DFT_r_v2_37_reset),
    .io_in_0_Re(DFT_r_v2_37_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_37_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_37_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_37_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_37_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_37_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_37_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_37_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_38 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_38_clock),
    .reset(DFT_r_v2_38_reset),
    .io_in_0_Re(DFT_r_v2_38_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_38_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_38_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_38_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_38_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_38_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_38_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_38_io_out_1_Im)
  );
  DFT_r_v2 DFT_r_v2_39 ( // @[FFTDesigns.scala 5100:30]
    .clock(DFT_r_v2_39_clock),
    .reset(DFT_r_v2_39_reset),
    .io_in_0_Re(DFT_r_v2_39_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_39_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_39_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_39_io_in_1_Im),
    .io_out_0_Re(DFT_r_v2_39_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_39_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_39_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_39_io_out_1_Im)
  );
  PermutationsWithStreaming PermutationsWithStreaming ( // @[FFTDesigns.scala 5107:30]
    .clock(PermutationsWithStreaming_clock),
    .reset(PermutationsWithStreaming_reset),
    .io_in_0_Re(PermutationsWithStreaming_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_io_in_15_Im),
    .io_in_en_0(PermutationsWithStreaming_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_io_in_en_4),
    .io_out_0_Re(PermutationsWithStreaming_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_io_out_15_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_1 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_1_clock),
    .reset(PermutationsWithStreaming_1_reset),
    .io_in_0_Re(PermutationsWithStreaming_1_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_1_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_1_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_1_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_1_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_1_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_1_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_1_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_1_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_1_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_1_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_1_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_1_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_1_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_1_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_1_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_1_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_1_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_1_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_1_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_1_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_1_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_1_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_1_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_1_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_1_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_1_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_1_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_1_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_1_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_1_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_1_io_in_15_Im),
    .io_in_en_0(PermutationsWithStreaming_1_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_1_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_1_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_1_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_1_io_in_en_4),
    .io_out_0_Re(PermutationsWithStreaming_1_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_1_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_1_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_1_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_1_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_1_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_1_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_1_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_1_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_1_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_1_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_1_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_1_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_1_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_1_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_1_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_1_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_1_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_1_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_1_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_1_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_1_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_1_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_1_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_1_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_1_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_1_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_1_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_1_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_1_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_1_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_1_io_out_15_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_2 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_2_clock),
    .reset(PermutationsWithStreaming_2_reset),
    .io_in_0_Re(PermutationsWithStreaming_2_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_2_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_2_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_2_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_2_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_2_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_2_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_2_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_2_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_2_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_2_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_2_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_2_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_2_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_2_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_2_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_2_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_2_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_2_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_2_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_2_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_2_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_2_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_2_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_2_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_2_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_2_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_2_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_2_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_2_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_2_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_2_io_in_15_Im),
    .io_in_en_0(PermutationsWithStreaming_2_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_2_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_2_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_2_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_2_io_in_en_4),
    .io_out_0_Re(PermutationsWithStreaming_2_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_2_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_2_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_2_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_2_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_2_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_2_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_2_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_2_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_2_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_2_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_2_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_2_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_2_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_2_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_2_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_2_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_2_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_2_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_2_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_2_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_2_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_2_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_2_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_2_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_2_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_2_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_2_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_2_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_2_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_2_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_2_io_out_15_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_3 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_3_clock),
    .reset(PermutationsWithStreaming_3_reset),
    .io_in_0_Re(PermutationsWithStreaming_3_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_3_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_3_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_3_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_3_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_3_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_3_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_3_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_3_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_3_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_3_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_3_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_3_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_3_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_3_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_3_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_3_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_3_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_3_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_3_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_3_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_3_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_3_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_3_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_3_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_3_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_3_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_3_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_3_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_3_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_3_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_3_io_in_15_Im),
    .io_in_en_0(PermutationsWithStreaming_3_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_3_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_3_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_3_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_3_io_in_en_4),
    .io_out_0_Re(PermutationsWithStreaming_3_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_3_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_3_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_3_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_3_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_3_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_3_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_3_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_3_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_3_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_3_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_3_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_3_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_3_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_3_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_3_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_3_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_3_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_3_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_3_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_3_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_3_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_3_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_3_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_3_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_3_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_3_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_3_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_3_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_3_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_3_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_3_io_out_15_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_4 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_4_clock),
    .reset(PermutationsWithStreaming_4_reset),
    .io_in_0_Re(PermutationsWithStreaming_4_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_4_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_4_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_4_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_4_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_4_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_4_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_4_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_4_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_4_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_4_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_4_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_4_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_4_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_4_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_4_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_4_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_4_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_4_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_4_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_4_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_4_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_4_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_4_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_4_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_4_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_4_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_4_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_4_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_4_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_4_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_4_io_in_15_Im),
    .io_in_en_0(PermutationsWithStreaming_4_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_4_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_4_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_4_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_4_io_in_en_4),
    .io_out_0_Re(PermutationsWithStreaming_4_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_4_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_4_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_4_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_4_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_4_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_4_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_4_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_4_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_4_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_4_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_4_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_4_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_4_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_4_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_4_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_4_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_4_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_4_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_4_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_4_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_4_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_4_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_4_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_4_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_4_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_4_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_4_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_4_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_4_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_4_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_4_io_out_15_Im)
  );
  PermutationsWithStreaming_1 PermutationsWithStreaming_5 ( // @[FFTDesigns.scala 5110:30]
    .clock(PermutationsWithStreaming_5_clock),
    .reset(PermutationsWithStreaming_5_reset),
    .io_in_0_Re(PermutationsWithStreaming_5_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_5_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_5_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_5_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_5_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_5_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_5_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_5_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_5_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_5_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_5_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_5_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_5_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_5_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_5_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_5_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_5_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_5_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_5_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_5_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_5_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_5_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_5_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_5_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_5_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_5_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_5_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_5_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_5_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_5_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_5_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_5_io_in_15_Im),
    .io_in_en_0(PermutationsWithStreaming_5_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_5_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_5_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_5_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_5_io_in_en_4),
    .io_out_0_Re(PermutationsWithStreaming_5_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_5_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_5_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_5_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_5_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_5_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_5_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_5_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_5_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_5_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_5_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_5_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_5_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_5_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_5_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_5_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_5_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_5_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_5_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_5_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_5_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_5_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_5_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_5_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_5_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_5_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_5_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_5_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_5_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_5_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_5_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_5_io_out_15_Im)
  );
  TwiddleFactorsStreamed TwiddleFactorsStreamed ( // @[FFTDesigns.scala 5115:28]
    .clock(TwiddleFactorsStreamed_clock),
    .reset(TwiddleFactorsStreamed_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_io_in_7_Im),
    .io_in_8_Re(TwiddleFactorsStreamed_io_in_8_Re),
    .io_in_8_Im(TwiddleFactorsStreamed_io_in_8_Im),
    .io_in_9_Re(TwiddleFactorsStreamed_io_in_9_Re),
    .io_in_9_Im(TwiddleFactorsStreamed_io_in_9_Im),
    .io_in_10_Re(TwiddleFactorsStreamed_io_in_10_Re),
    .io_in_10_Im(TwiddleFactorsStreamed_io_in_10_Im),
    .io_in_11_Re(TwiddleFactorsStreamed_io_in_11_Re),
    .io_in_11_Im(TwiddleFactorsStreamed_io_in_11_Im),
    .io_in_12_Re(TwiddleFactorsStreamed_io_in_12_Re),
    .io_in_12_Im(TwiddleFactorsStreamed_io_in_12_Im),
    .io_in_13_Re(TwiddleFactorsStreamed_io_in_13_Re),
    .io_in_13_Im(TwiddleFactorsStreamed_io_in_13_Im),
    .io_in_14_Re(TwiddleFactorsStreamed_io_in_14_Re),
    .io_in_14_Im(TwiddleFactorsStreamed_io_in_14_Im),
    .io_in_15_Re(TwiddleFactorsStreamed_io_in_15_Re),
    .io_in_15_Im(TwiddleFactorsStreamed_io_in_15_Im),
    .io_in_en_0(TwiddleFactorsStreamed_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_io_out_7_Im),
    .io_out_8_Re(TwiddleFactorsStreamed_io_out_8_Re),
    .io_out_8_Im(TwiddleFactorsStreamed_io_out_8_Im),
    .io_out_9_Re(TwiddleFactorsStreamed_io_out_9_Re),
    .io_out_9_Im(TwiddleFactorsStreamed_io_out_9_Im),
    .io_out_10_Re(TwiddleFactorsStreamed_io_out_10_Re),
    .io_out_10_Im(TwiddleFactorsStreamed_io_out_10_Im),
    .io_out_11_Re(TwiddleFactorsStreamed_io_out_11_Re),
    .io_out_11_Im(TwiddleFactorsStreamed_io_out_11_Im),
    .io_out_12_Re(TwiddleFactorsStreamed_io_out_12_Re),
    .io_out_12_Im(TwiddleFactorsStreamed_io_out_12_Im),
    .io_out_13_Re(TwiddleFactorsStreamed_io_out_13_Re),
    .io_out_13_Im(TwiddleFactorsStreamed_io_out_13_Im),
    .io_out_14_Re(TwiddleFactorsStreamed_io_out_14_Re),
    .io_out_14_Im(TwiddleFactorsStreamed_io_out_14_Im),
    .io_out_15_Re(TwiddleFactorsStreamed_io_out_15_Re),
    .io_out_15_Im(TwiddleFactorsStreamed_io_out_15_Im)
  );
  TwiddleFactorsStreamed_1 TwiddleFactorsStreamed_1 ( // @[FFTDesigns.scala 5115:28]
    .clock(TwiddleFactorsStreamed_1_clock),
    .reset(TwiddleFactorsStreamed_1_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_1_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_1_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_1_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_1_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_1_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_1_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_1_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_1_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_1_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_1_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_1_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_1_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_1_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_1_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_1_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_1_io_in_7_Im),
    .io_in_8_Re(TwiddleFactorsStreamed_1_io_in_8_Re),
    .io_in_8_Im(TwiddleFactorsStreamed_1_io_in_8_Im),
    .io_in_9_Re(TwiddleFactorsStreamed_1_io_in_9_Re),
    .io_in_9_Im(TwiddleFactorsStreamed_1_io_in_9_Im),
    .io_in_10_Re(TwiddleFactorsStreamed_1_io_in_10_Re),
    .io_in_10_Im(TwiddleFactorsStreamed_1_io_in_10_Im),
    .io_in_11_Re(TwiddleFactorsStreamed_1_io_in_11_Re),
    .io_in_11_Im(TwiddleFactorsStreamed_1_io_in_11_Im),
    .io_in_12_Re(TwiddleFactorsStreamed_1_io_in_12_Re),
    .io_in_12_Im(TwiddleFactorsStreamed_1_io_in_12_Im),
    .io_in_13_Re(TwiddleFactorsStreamed_1_io_in_13_Re),
    .io_in_13_Im(TwiddleFactorsStreamed_1_io_in_13_Im),
    .io_in_14_Re(TwiddleFactorsStreamed_1_io_in_14_Re),
    .io_in_14_Im(TwiddleFactorsStreamed_1_io_in_14_Im),
    .io_in_15_Re(TwiddleFactorsStreamed_1_io_in_15_Re),
    .io_in_15_Im(TwiddleFactorsStreamed_1_io_in_15_Im),
    .io_in_en_0(TwiddleFactorsStreamed_1_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_1_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_1_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_1_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_1_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_1_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_1_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_1_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_1_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_1_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_1_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_1_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_1_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_1_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_1_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_1_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_1_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_1_io_out_7_Im),
    .io_out_8_Re(TwiddleFactorsStreamed_1_io_out_8_Re),
    .io_out_8_Im(TwiddleFactorsStreamed_1_io_out_8_Im),
    .io_out_9_Re(TwiddleFactorsStreamed_1_io_out_9_Re),
    .io_out_9_Im(TwiddleFactorsStreamed_1_io_out_9_Im),
    .io_out_10_Re(TwiddleFactorsStreamed_1_io_out_10_Re),
    .io_out_10_Im(TwiddleFactorsStreamed_1_io_out_10_Im),
    .io_out_11_Re(TwiddleFactorsStreamed_1_io_out_11_Re),
    .io_out_11_Im(TwiddleFactorsStreamed_1_io_out_11_Im),
    .io_out_12_Re(TwiddleFactorsStreamed_1_io_out_12_Re),
    .io_out_12_Im(TwiddleFactorsStreamed_1_io_out_12_Im),
    .io_out_13_Re(TwiddleFactorsStreamed_1_io_out_13_Re),
    .io_out_13_Im(TwiddleFactorsStreamed_1_io_out_13_Im),
    .io_out_14_Re(TwiddleFactorsStreamed_1_io_out_14_Re),
    .io_out_14_Im(TwiddleFactorsStreamed_1_io_out_14_Im),
    .io_out_15_Re(TwiddleFactorsStreamed_1_io_out_15_Re),
    .io_out_15_Im(TwiddleFactorsStreamed_1_io_out_15_Im)
  );
  TwiddleFactorsStreamed_2 TwiddleFactorsStreamed_2 ( // @[FFTDesigns.scala 5115:28]
    .clock(TwiddleFactorsStreamed_2_clock),
    .reset(TwiddleFactorsStreamed_2_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_2_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_2_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_2_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_2_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_2_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_2_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_2_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_2_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_2_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_2_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_2_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_2_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_2_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_2_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_2_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_2_io_in_7_Im),
    .io_in_8_Re(TwiddleFactorsStreamed_2_io_in_8_Re),
    .io_in_8_Im(TwiddleFactorsStreamed_2_io_in_8_Im),
    .io_in_9_Re(TwiddleFactorsStreamed_2_io_in_9_Re),
    .io_in_9_Im(TwiddleFactorsStreamed_2_io_in_9_Im),
    .io_in_10_Re(TwiddleFactorsStreamed_2_io_in_10_Re),
    .io_in_10_Im(TwiddleFactorsStreamed_2_io_in_10_Im),
    .io_in_11_Re(TwiddleFactorsStreamed_2_io_in_11_Re),
    .io_in_11_Im(TwiddleFactorsStreamed_2_io_in_11_Im),
    .io_in_12_Re(TwiddleFactorsStreamed_2_io_in_12_Re),
    .io_in_12_Im(TwiddleFactorsStreamed_2_io_in_12_Im),
    .io_in_13_Re(TwiddleFactorsStreamed_2_io_in_13_Re),
    .io_in_13_Im(TwiddleFactorsStreamed_2_io_in_13_Im),
    .io_in_14_Re(TwiddleFactorsStreamed_2_io_in_14_Re),
    .io_in_14_Im(TwiddleFactorsStreamed_2_io_in_14_Im),
    .io_in_15_Re(TwiddleFactorsStreamed_2_io_in_15_Re),
    .io_in_15_Im(TwiddleFactorsStreamed_2_io_in_15_Im),
    .io_in_en_0(TwiddleFactorsStreamed_2_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_2_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_2_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_2_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_2_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_2_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_2_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_2_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_2_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_2_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_2_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_2_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_2_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_2_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_2_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_2_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_2_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_2_io_out_7_Im),
    .io_out_8_Re(TwiddleFactorsStreamed_2_io_out_8_Re),
    .io_out_8_Im(TwiddleFactorsStreamed_2_io_out_8_Im),
    .io_out_9_Re(TwiddleFactorsStreamed_2_io_out_9_Re),
    .io_out_9_Im(TwiddleFactorsStreamed_2_io_out_9_Im),
    .io_out_10_Re(TwiddleFactorsStreamed_2_io_out_10_Re),
    .io_out_10_Im(TwiddleFactorsStreamed_2_io_out_10_Im),
    .io_out_11_Re(TwiddleFactorsStreamed_2_io_out_11_Re),
    .io_out_11_Im(TwiddleFactorsStreamed_2_io_out_11_Im),
    .io_out_12_Re(TwiddleFactorsStreamed_2_io_out_12_Re),
    .io_out_12_Im(TwiddleFactorsStreamed_2_io_out_12_Im),
    .io_out_13_Re(TwiddleFactorsStreamed_2_io_out_13_Re),
    .io_out_13_Im(TwiddleFactorsStreamed_2_io_out_13_Im),
    .io_out_14_Re(TwiddleFactorsStreamed_2_io_out_14_Re),
    .io_out_14_Im(TwiddleFactorsStreamed_2_io_out_14_Im),
    .io_out_15_Re(TwiddleFactorsStreamed_2_io_out_15_Re),
    .io_out_15_Im(TwiddleFactorsStreamed_2_io_out_15_Im)
  );
  TwiddleFactorsStreamed_3 TwiddleFactorsStreamed_3 ( // @[FFTDesigns.scala 5115:28]
    .clock(TwiddleFactorsStreamed_3_clock),
    .reset(TwiddleFactorsStreamed_3_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_3_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_3_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_3_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_3_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_3_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_3_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_3_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_3_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_3_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_3_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_3_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_3_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_3_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_3_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_3_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_3_io_in_7_Im),
    .io_in_8_Re(TwiddleFactorsStreamed_3_io_in_8_Re),
    .io_in_8_Im(TwiddleFactorsStreamed_3_io_in_8_Im),
    .io_in_9_Re(TwiddleFactorsStreamed_3_io_in_9_Re),
    .io_in_9_Im(TwiddleFactorsStreamed_3_io_in_9_Im),
    .io_in_10_Re(TwiddleFactorsStreamed_3_io_in_10_Re),
    .io_in_10_Im(TwiddleFactorsStreamed_3_io_in_10_Im),
    .io_in_11_Re(TwiddleFactorsStreamed_3_io_in_11_Re),
    .io_in_11_Im(TwiddleFactorsStreamed_3_io_in_11_Im),
    .io_in_12_Re(TwiddleFactorsStreamed_3_io_in_12_Re),
    .io_in_12_Im(TwiddleFactorsStreamed_3_io_in_12_Im),
    .io_in_13_Re(TwiddleFactorsStreamed_3_io_in_13_Re),
    .io_in_13_Im(TwiddleFactorsStreamed_3_io_in_13_Im),
    .io_in_14_Re(TwiddleFactorsStreamed_3_io_in_14_Re),
    .io_in_14_Im(TwiddleFactorsStreamed_3_io_in_14_Im),
    .io_in_15_Re(TwiddleFactorsStreamed_3_io_in_15_Re),
    .io_in_15_Im(TwiddleFactorsStreamed_3_io_in_15_Im),
    .io_in_en_0(TwiddleFactorsStreamed_3_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_3_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_3_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_3_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_3_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_3_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_3_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_3_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_3_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_3_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_3_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_3_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_3_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_3_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_3_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_3_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_3_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_3_io_out_7_Im),
    .io_out_8_Re(TwiddleFactorsStreamed_3_io_out_8_Re),
    .io_out_8_Im(TwiddleFactorsStreamed_3_io_out_8_Im),
    .io_out_9_Re(TwiddleFactorsStreamed_3_io_out_9_Re),
    .io_out_9_Im(TwiddleFactorsStreamed_3_io_out_9_Im),
    .io_out_10_Re(TwiddleFactorsStreamed_3_io_out_10_Re),
    .io_out_10_Im(TwiddleFactorsStreamed_3_io_out_10_Im),
    .io_out_11_Re(TwiddleFactorsStreamed_3_io_out_11_Re),
    .io_out_11_Im(TwiddleFactorsStreamed_3_io_out_11_Im),
    .io_out_12_Re(TwiddleFactorsStreamed_3_io_out_12_Re),
    .io_out_12_Im(TwiddleFactorsStreamed_3_io_out_12_Im),
    .io_out_13_Re(TwiddleFactorsStreamed_3_io_out_13_Re),
    .io_out_13_Im(TwiddleFactorsStreamed_3_io_out_13_Im),
    .io_out_14_Re(TwiddleFactorsStreamed_3_io_out_14_Re),
    .io_out_14_Im(TwiddleFactorsStreamed_3_io_out_14_Im),
    .io_out_15_Re(TwiddleFactorsStreamed_3_io_out_15_Re),
    .io_out_15_Im(TwiddleFactorsStreamed_3_io_out_15_Im)
  );
  assign io_out_0_Re = PermutationsWithStreaming_5_io_out_0_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_0_Im = PermutationsWithStreaming_5_io_out_0_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_1_Re = PermutationsWithStreaming_5_io_out_1_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_1_Im = PermutationsWithStreaming_5_io_out_1_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_2_Re = PermutationsWithStreaming_5_io_out_2_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_2_Im = PermutationsWithStreaming_5_io_out_2_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_3_Re = PermutationsWithStreaming_5_io_out_3_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_3_Im = PermutationsWithStreaming_5_io_out_3_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_4_Re = PermutationsWithStreaming_5_io_out_4_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_4_Im = PermutationsWithStreaming_5_io_out_4_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_5_Re = PermutationsWithStreaming_5_io_out_5_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_5_Im = PermutationsWithStreaming_5_io_out_5_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_6_Re = PermutationsWithStreaming_5_io_out_6_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_6_Im = PermutationsWithStreaming_5_io_out_6_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_7_Re = PermutationsWithStreaming_5_io_out_7_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_7_Im = PermutationsWithStreaming_5_io_out_7_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_8_Re = PermutationsWithStreaming_5_io_out_8_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_8_Im = PermutationsWithStreaming_5_io_out_8_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_9_Re = PermutationsWithStreaming_5_io_out_9_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_9_Im = PermutationsWithStreaming_5_io_out_9_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_10_Re = PermutationsWithStreaming_5_io_out_10_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_10_Im = PermutationsWithStreaming_5_io_out_10_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_11_Re = PermutationsWithStreaming_5_io_out_11_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_11_Im = PermutationsWithStreaming_5_io_out_11_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_12_Re = PermutationsWithStreaming_5_io_out_12_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_12_Im = PermutationsWithStreaming_5_io_out_12_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_13_Re = PermutationsWithStreaming_5_io_out_13_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_13_Im = PermutationsWithStreaming_5_io_out_13_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_14_Re = PermutationsWithStreaming_5_io_out_14_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_14_Im = PermutationsWithStreaming_5_io_out_14_Im; // @[FFTDesigns.scala 5201:12]
  assign io_out_15_Re = PermutationsWithStreaming_5_io_out_15_Re; // @[FFTDesigns.scala 5201:12]
  assign io_out_15_Im = PermutationsWithStreaming_5_io_out_15_Im; // @[FFTDesigns.scala 5201:12]
  assign DFT_r_v2_clock = clock;
  assign DFT_r_v2_reset = reset;
  assign DFT_r_v2_io_in_0_Re = PermutationsWithStreaming_io_out_0_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_io_in_0_Im = PermutationsWithStreaming_io_out_0_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_io_in_1_Re = PermutationsWithStreaming_io_out_1_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_io_in_1_Im = PermutationsWithStreaming_io_out_1_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_1_clock = clock;
  assign DFT_r_v2_1_reset = reset;
  assign DFT_r_v2_1_io_in_0_Re = PermutationsWithStreaming_io_out_2_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_1_io_in_0_Im = PermutationsWithStreaming_io_out_2_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_1_io_in_1_Re = PermutationsWithStreaming_io_out_3_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_1_io_in_1_Im = PermutationsWithStreaming_io_out_3_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_2_clock = clock;
  assign DFT_r_v2_2_reset = reset;
  assign DFT_r_v2_2_io_in_0_Re = PermutationsWithStreaming_io_out_4_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_2_io_in_0_Im = PermutationsWithStreaming_io_out_4_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_2_io_in_1_Re = PermutationsWithStreaming_io_out_5_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_2_io_in_1_Im = PermutationsWithStreaming_io_out_5_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_3_clock = clock;
  assign DFT_r_v2_3_reset = reset;
  assign DFT_r_v2_3_io_in_0_Re = PermutationsWithStreaming_io_out_6_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_3_io_in_0_Im = PermutationsWithStreaming_io_out_6_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_3_io_in_1_Re = PermutationsWithStreaming_io_out_7_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_3_io_in_1_Im = PermutationsWithStreaming_io_out_7_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_4_clock = clock;
  assign DFT_r_v2_4_reset = reset;
  assign DFT_r_v2_4_io_in_0_Re = PermutationsWithStreaming_io_out_8_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_4_io_in_0_Im = PermutationsWithStreaming_io_out_8_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_4_io_in_1_Re = PermutationsWithStreaming_io_out_9_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_4_io_in_1_Im = PermutationsWithStreaming_io_out_9_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_5_clock = clock;
  assign DFT_r_v2_5_reset = reset;
  assign DFT_r_v2_5_io_in_0_Re = PermutationsWithStreaming_io_out_10_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_5_io_in_0_Im = PermutationsWithStreaming_io_out_10_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_5_io_in_1_Re = PermutationsWithStreaming_io_out_11_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_5_io_in_1_Im = PermutationsWithStreaming_io_out_11_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_6_clock = clock;
  assign DFT_r_v2_6_reset = reset;
  assign DFT_r_v2_6_io_in_0_Re = PermutationsWithStreaming_io_out_12_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_6_io_in_0_Im = PermutationsWithStreaming_io_out_12_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_6_io_in_1_Re = PermutationsWithStreaming_io_out_13_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_6_io_in_1_Im = PermutationsWithStreaming_io_out_13_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_7_clock = clock;
  assign DFT_r_v2_7_reset = reset;
  assign DFT_r_v2_7_io_in_0_Re = PermutationsWithStreaming_io_out_14_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_7_io_in_0_Im = PermutationsWithStreaming_io_out_14_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_7_io_in_1_Re = PermutationsWithStreaming_io_out_15_Re; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_7_io_in_1_Im = PermutationsWithStreaming_io_out_15_Im; // @[FFTDesigns.scala 5156:41]
  assign DFT_r_v2_8_clock = clock;
  assign DFT_r_v2_8_reset = reset;
  assign DFT_r_v2_8_io_in_0_Re = TwiddleFactorsStreamed_io_out_0_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_8_io_in_0_Im = TwiddleFactorsStreamed_io_out_0_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_8_io_in_1_Re = TwiddleFactorsStreamed_io_out_1_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_8_io_in_1_Im = TwiddleFactorsStreamed_io_out_1_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_9_clock = clock;
  assign DFT_r_v2_9_reset = reset;
  assign DFT_r_v2_9_io_in_0_Re = TwiddleFactorsStreamed_io_out_2_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_9_io_in_0_Im = TwiddleFactorsStreamed_io_out_2_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_9_io_in_1_Re = TwiddleFactorsStreamed_io_out_3_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_9_io_in_1_Im = TwiddleFactorsStreamed_io_out_3_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_10_clock = clock;
  assign DFT_r_v2_10_reset = reset;
  assign DFT_r_v2_10_io_in_0_Re = TwiddleFactorsStreamed_io_out_4_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_10_io_in_0_Im = TwiddleFactorsStreamed_io_out_4_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_10_io_in_1_Re = TwiddleFactorsStreamed_io_out_5_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_10_io_in_1_Im = TwiddleFactorsStreamed_io_out_5_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_11_clock = clock;
  assign DFT_r_v2_11_reset = reset;
  assign DFT_r_v2_11_io_in_0_Re = TwiddleFactorsStreamed_io_out_6_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_11_io_in_0_Im = TwiddleFactorsStreamed_io_out_6_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_11_io_in_1_Re = TwiddleFactorsStreamed_io_out_7_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_11_io_in_1_Im = TwiddleFactorsStreamed_io_out_7_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_12_clock = clock;
  assign DFT_r_v2_12_reset = reset;
  assign DFT_r_v2_12_io_in_0_Re = TwiddleFactorsStreamed_io_out_8_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_12_io_in_0_Im = TwiddleFactorsStreamed_io_out_8_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_12_io_in_1_Re = TwiddleFactorsStreamed_io_out_9_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_12_io_in_1_Im = TwiddleFactorsStreamed_io_out_9_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_13_clock = clock;
  assign DFT_r_v2_13_reset = reset;
  assign DFT_r_v2_13_io_in_0_Re = TwiddleFactorsStreamed_io_out_10_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_13_io_in_0_Im = TwiddleFactorsStreamed_io_out_10_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_13_io_in_1_Re = TwiddleFactorsStreamed_io_out_11_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_13_io_in_1_Im = TwiddleFactorsStreamed_io_out_11_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_14_clock = clock;
  assign DFT_r_v2_14_reset = reset;
  assign DFT_r_v2_14_io_in_0_Re = TwiddleFactorsStreamed_io_out_12_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_14_io_in_0_Im = TwiddleFactorsStreamed_io_out_12_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_14_io_in_1_Re = TwiddleFactorsStreamed_io_out_13_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_14_io_in_1_Im = TwiddleFactorsStreamed_io_out_13_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_15_clock = clock;
  assign DFT_r_v2_15_reset = reset;
  assign DFT_r_v2_15_io_in_0_Re = TwiddleFactorsStreamed_io_out_14_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_15_io_in_0_Im = TwiddleFactorsStreamed_io_out_14_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_15_io_in_1_Re = TwiddleFactorsStreamed_io_out_15_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_15_io_in_1_Im = TwiddleFactorsStreamed_io_out_15_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_16_clock = clock;
  assign DFT_r_v2_16_reset = reset;
  assign DFT_r_v2_16_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_0_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_16_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_0_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_16_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_1_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_16_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_1_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_17_clock = clock;
  assign DFT_r_v2_17_reset = reset;
  assign DFT_r_v2_17_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_2_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_17_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_2_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_17_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_3_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_17_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_3_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_18_clock = clock;
  assign DFT_r_v2_18_reset = reset;
  assign DFT_r_v2_18_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_4_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_18_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_4_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_18_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_5_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_18_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_5_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_19_clock = clock;
  assign DFT_r_v2_19_reset = reset;
  assign DFT_r_v2_19_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_6_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_19_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_6_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_19_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_7_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_19_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_7_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_20_clock = clock;
  assign DFT_r_v2_20_reset = reset;
  assign DFT_r_v2_20_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_8_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_20_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_8_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_20_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_9_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_20_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_9_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_21_clock = clock;
  assign DFT_r_v2_21_reset = reset;
  assign DFT_r_v2_21_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_10_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_21_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_10_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_21_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_11_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_21_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_11_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_22_clock = clock;
  assign DFT_r_v2_22_reset = reset;
  assign DFT_r_v2_22_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_12_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_22_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_12_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_22_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_13_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_22_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_13_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_23_clock = clock;
  assign DFT_r_v2_23_reset = reset;
  assign DFT_r_v2_23_io_in_0_Re = TwiddleFactorsStreamed_1_io_out_14_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_23_io_in_0_Im = TwiddleFactorsStreamed_1_io_out_14_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_23_io_in_1_Re = TwiddleFactorsStreamed_1_io_out_15_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_23_io_in_1_Im = TwiddleFactorsStreamed_1_io_out_15_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_24_clock = clock;
  assign DFT_r_v2_24_reset = reset;
  assign DFT_r_v2_24_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_0_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_24_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_0_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_24_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_1_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_24_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_1_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_25_clock = clock;
  assign DFT_r_v2_25_reset = reset;
  assign DFT_r_v2_25_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_2_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_25_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_2_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_25_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_3_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_25_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_3_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_26_clock = clock;
  assign DFT_r_v2_26_reset = reset;
  assign DFT_r_v2_26_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_4_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_26_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_4_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_26_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_5_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_26_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_5_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_27_clock = clock;
  assign DFT_r_v2_27_reset = reset;
  assign DFT_r_v2_27_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_6_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_27_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_6_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_27_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_7_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_27_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_7_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_28_clock = clock;
  assign DFT_r_v2_28_reset = reset;
  assign DFT_r_v2_28_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_8_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_28_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_8_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_28_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_9_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_28_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_9_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_29_clock = clock;
  assign DFT_r_v2_29_reset = reset;
  assign DFT_r_v2_29_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_10_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_29_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_10_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_29_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_11_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_29_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_11_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_30_clock = clock;
  assign DFT_r_v2_30_reset = reset;
  assign DFT_r_v2_30_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_12_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_30_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_12_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_30_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_13_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_30_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_13_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_31_clock = clock;
  assign DFT_r_v2_31_reset = reset;
  assign DFT_r_v2_31_io_in_0_Re = TwiddleFactorsStreamed_2_io_out_14_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_31_io_in_0_Im = TwiddleFactorsStreamed_2_io_out_14_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_31_io_in_1_Re = TwiddleFactorsStreamed_2_io_out_15_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_31_io_in_1_Im = TwiddleFactorsStreamed_2_io_out_15_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_32_clock = clock;
  assign DFT_r_v2_32_reset = reset;
  assign DFT_r_v2_32_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_0_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_32_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_0_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_32_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_1_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_32_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_1_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_33_clock = clock;
  assign DFT_r_v2_33_reset = reset;
  assign DFT_r_v2_33_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_2_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_33_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_2_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_33_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_3_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_33_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_3_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_34_clock = clock;
  assign DFT_r_v2_34_reset = reset;
  assign DFT_r_v2_34_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_4_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_34_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_4_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_34_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_5_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_34_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_5_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_35_clock = clock;
  assign DFT_r_v2_35_reset = reset;
  assign DFT_r_v2_35_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_6_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_35_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_6_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_35_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_7_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_35_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_7_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_36_clock = clock;
  assign DFT_r_v2_36_reset = reset;
  assign DFT_r_v2_36_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_8_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_36_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_8_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_36_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_9_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_36_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_9_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_37_clock = clock;
  assign DFT_r_v2_37_reset = reset;
  assign DFT_r_v2_37_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_10_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_37_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_10_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_37_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_11_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_37_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_11_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_38_clock = clock;
  assign DFT_r_v2_38_reset = reset;
  assign DFT_r_v2_38_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_12_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_38_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_12_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_38_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_13_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_38_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_13_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_39_clock = clock;
  assign DFT_r_v2_39_reset = reset;
  assign DFT_r_v2_39_io_in_0_Re = TwiddleFactorsStreamed_3_io_out_14_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_39_io_in_0_Im = TwiddleFactorsStreamed_3_io_out_14_Im; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_39_io_in_1_Re = TwiddleFactorsStreamed_3_io_out_15_Re; // @[FFTDesigns.scala 5163:41]
  assign DFT_r_v2_39_io_in_1_Im = TwiddleFactorsStreamed_3_io_out_15_Im; // @[FFTDesigns.scala 5163:41]
  assign PermutationsWithStreaming_clock = clock;
  assign PermutationsWithStreaming_reset = reset;
  assign PermutationsWithStreaming_io_in_0_Re = io_in_ready ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_0_Im = io_in_ready ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_1_Re = io_in_ready ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_1_Im = io_in_ready ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_2_Re = io_in_ready ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_2_Im = io_in_ready ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_3_Re = io_in_ready ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_3_Im = io_in_ready ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_4_Re = io_in_ready ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_4_Im = io_in_ready ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_5_Re = io_in_ready ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_5_Im = io_in_ready ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_6_Re = io_in_ready ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_6_Im = io_in_ready ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_7_Re = io_in_ready ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_7_Im = io_in_ready ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_8_Re = io_in_ready ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_8_Im = io_in_ready ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_9_Re = io_in_ready ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_9_Im = io_in_ready ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_10_Re = io_in_ready ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_10_Im = io_in_ready ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_11_Re = io_in_ready ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_11_Im = io_in_ready ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_12_Re = io_in_ready ? io_in_12_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_12_Im = io_in_ready ? io_in_12_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_13_Re = io_in_ready ? io_in_13_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_13_Im = io_in_ready ? io_in_13_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_14_Re = io_in_ready ? io_in_14_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_14_Im = io_in_ready ? io_in_14_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_15_Re = io_in_ready ? io_in_15_Re : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_15_Im = io_in_ready ? io_in_15_Im : 32'h0; // @[FFTDesigns.scala 5124:30 5125:34 5128:39]
  assign PermutationsWithStreaming_io_in_en_0 = io_in_ready; // @[FFTDesigns.scala 5123:38]
  assign PermutationsWithStreaming_io_in_en_1 = Perm_regdelays_0_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_2 = Perm_regdelays_0_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_3 = Perm_regdelays_0_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_io_in_en_4 = Perm_regdelays_0_3; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_1_clock = clock;
  assign PermutationsWithStreaming_1_reset = reset;
  assign PermutationsWithStreaming_1_io_in_0_Re = DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_0_Im = DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_1_Re = DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_1_Im = DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_2_Re = DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_2_Im = DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_3_Re = DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_3_Im = DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_4_Re = DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_4_Im = DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_5_Re = DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_5_Im = DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_6_Re = DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_6_Im = DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_7_Re = DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_7_Im = DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_8_Re = DFT_r_v2_4_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_8_Im = DFT_r_v2_4_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_9_Re = DFT_r_v2_4_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_9_Im = DFT_r_v2_4_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_10_Re = DFT_r_v2_5_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_10_Im = DFT_r_v2_5_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_11_Re = DFT_r_v2_5_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_11_Im = DFT_r_v2_5_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_12_Re = DFT_r_v2_6_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_12_Im = DFT_r_v2_6_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_13_Re = DFT_r_v2_6_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_13_Im = DFT_r_v2_6_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_14_Re = DFT_r_v2_7_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_14_Im = DFT_r_v2_7_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_15_Re = DFT_r_v2_7_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_15_Im = DFT_r_v2_7_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_1_io_in_en_0 = DFT_regdelays_0_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_1_io_in_en_1 = Perm_regdelays_1_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_2 = Perm_regdelays_1_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_3 = Perm_regdelays_1_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_1_io_in_en_4 = Perm_regdelays_1_3; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_2_clock = clock;
  assign PermutationsWithStreaming_2_reset = reset;
  assign PermutationsWithStreaming_2_io_in_0_Re = DFT_r_v2_8_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_0_Im = DFT_r_v2_8_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_1_Re = DFT_r_v2_8_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_1_Im = DFT_r_v2_8_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_2_Re = DFT_r_v2_9_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_2_Im = DFT_r_v2_9_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_3_Re = DFT_r_v2_9_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_3_Im = DFT_r_v2_9_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_4_Re = DFT_r_v2_10_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_4_Im = DFT_r_v2_10_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_5_Re = DFT_r_v2_10_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_5_Im = DFT_r_v2_10_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_6_Re = DFT_r_v2_11_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_6_Im = DFT_r_v2_11_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_7_Re = DFT_r_v2_11_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_7_Im = DFT_r_v2_11_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_8_Re = DFT_r_v2_12_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_8_Im = DFT_r_v2_12_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_9_Re = DFT_r_v2_12_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_9_Im = DFT_r_v2_12_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_10_Re = DFT_r_v2_13_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_10_Im = DFT_r_v2_13_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_11_Re = DFT_r_v2_13_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_11_Im = DFT_r_v2_13_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_12_Re = DFT_r_v2_14_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_12_Im = DFT_r_v2_14_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_13_Re = DFT_r_v2_14_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_13_Im = DFT_r_v2_14_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_14_Re = DFT_r_v2_15_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_14_Im = DFT_r_v2_15_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_15_Re = DFT_r_v2_15_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_15_Im = DFT_r_v2_15_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_2_io_in_en_0 = DFT_regdelays_1_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_2_io_in_en_1 = Perm_regdelays_2_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_2 = Perm_regdelays_2_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_3 = Perm_regdelays_2_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_2_io_in_en_4 = Perm_regdelays_2_3; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_3_clock = clock;
  assign PermutationsWithStreaming_3_reset = reset;
  assign PermutationsWithStreaming_3_io_in_0_Re = DFT_r_v2_16_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_0_Im = DFT_r_v2_16_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_1_Re = DFT_r_v2_16_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_1_Im = DFT_r_v2_16_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_2_Re = DFT_r_v2_17_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_2_Im = DFT_r_v2_17_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_3_Re = DFT_r_v2_17_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_3_Im = DFT_r_v2_17_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_4_Re = DFT_r_v2_18_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_4_Im = DFT_r_v2_18_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_5_Re = DFT_r_v2_18_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_5_Im = DFT_r_v2_18_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_6_Re = DFT_r_v2_19_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_6_Im = DFT_r_v2_19_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_7_Re = DFT_r_v2_19_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_7_Im = DFT_r_v2_19_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_8_Re = DFT_r_v2_20_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_8_Im = DFT_r_v2_20_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_9_Re = DFT_r_v2_20_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_9_Im = DFT_r_v2_20_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_10_Re = DFT_r_v2_21_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_10_Im = DFT_r_v2_21_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_11_Re = DFT_r_v2_21_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_11_Im = DFT_r_v2_21_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_12_Re = DFT_r_v2_22_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_12_Im = DFT_r_v2_22_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_13_Re = DFT_r_v2_22_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_13_Im = DFT_r_v2_22_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_14_Re = DFT_r_v2_23_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_14_Im = DFT_r_v2_23_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_15_Re = DFT_r_v2_23_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_15_Im = DFT_r_v2_23_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_3_io_in_en_0 = DFT_regdelays_2_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_3_io_in_en_1 = Perm_regdelays_3_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_2 = Perm_regdelays_3_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_3 = Perm_regdelays_3_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_3_io_in_en_4 = Perm_regdelays_3_3; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_4_clock = clock;
  assign PermutationsWithStreaming_4_reset = reset;
  assign PermutationsWithStreaming_4_io_in_0_Re = DFT_r_v2_24_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_0_Im = DFT_r_v2_24_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_1_Re = DFT_r_v2_24_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_1_Im = DFT_r_v2_24_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_2_Re = DFT_r_v2_25_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_2_Im = DFT_r_v2_25_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_3_Re = DFT_r_v2_25_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_3_Im = DFT_r_v2_25_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_4_Re = DFT_r_v2_26_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_4_Im = DFT_r_v2_26_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_5_Re = DFT_r_v2_26_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_5_Im = DFT_r_v2_26_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_6_Re = DFT_r_v2_27_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_6_Im = DFT_r_v2_27_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_7_Re = DFT_r_v2_27_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_7_Im = DFT_r_v2_27_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_8_Re = DFT_r_v2_28_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_8_Im = DFT_r_v2_28_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_9_Re = DFT_r_v2_28_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_9_Im = DFT_r_v2_28_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_10_Re = DFT_r_v2_29_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_10_Im = DFT_r_v2_29_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_11_Re = DFT_r_v2_29_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_11_Im = DFT_r_v2_29_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_12_Re = DFT_r_v2_30_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_12_Im = DFT_r_v2_30_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_13_Re = DFT_r_v2_30_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_13_Im = DFT_r_v2_30_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_14_Re = DFT_r_v2_31_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_14_Im = DFT_r_v2_31_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_15_Re = DFT_r_v2_31_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_15_Im = DFT_r_v2_31_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_4_io_in_en_0 = DFT_regdelays_3_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_4_io_in_en_1 = Perm_regdelays_4_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_2 = Perm_regdelays_4_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_3 = Perm_regdelays_4_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_4_io_in_en_4 = Perm_regdelays_4_3; // @[FFTDesigns.scala 5144:44]
  assign PermutationsWithStreaming_5_clock = clock;
  assign PermutationsWithStreaming_5_reset = reset;
  assign PermutationsWithStreaming_5_io_in_0_Re = DFT_r_v2_32_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_0_Im = DFT_r_v2_32_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_1_Re = DFT_r_v2_32_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_1_Im = DFT_r_v2_32_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_2_Re = DFT_r_v2_33_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_2_Im = DFT_r_v2_33_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_3_Re = DFT_r_v2_33_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_3_Im = DFT_r_v2_33_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_4_Re = DFT_r_v2_34_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_4_Im = DFT_r_v2_34_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_5_Re = DFT_r_v2_34_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_5_Im = DFT_r_v2_34_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_6_Re = DFT_r_v2_35_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_6_Im = DFT_r_v2_35_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_7_Re = DFT_r_v2_35_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_7_Im = DFT_r_v2_35_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_8_Re = DFT_r_v2_36_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_8_Im = DFT_r_v2_36_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_9_Re = DFT_r_v2_36_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_9_Im = DFT_r_v2_36_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_10_Re = DFT_r_v2_37_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_10_Im = DFT_r_v2_37_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_11_Re = DFT_r_v2_37_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_11_Im = DFT_r_v2_37_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_12_Re = DFT_r_v2_38_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_12_Im = DFT_r_v2_38_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_13_Re = DFT_r_v2_38_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_13_Im = DFT_r_v2_38_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_14_Re = DFT_r_v2_39_io_out_0_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_14_Im = DFT_r_v2_39_io_out_0_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_15_Re = DFT_r_v2_39_io_out_1_Re; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_15_Im = DFT_r_v2_39_io_out_1_Im; // @[FFTDesigns.scala 5136:45]
  assign PermutationsWithStreaming_5_io_in_en_0 = DFT_regdelays_4_0; // @[FFTDesigns.scala 5133:38]
  assign PermutationsWithStreaming_5_io_in_en_1 = Perm_regdelays_5_0; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_2 = Perm_regdelays_5_1; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_3 = Perm_regdelays_5_2; // @[FFTDesigns.scala 5142:36]
  assign PermutationsWithStreaming_5_io_in_en_4 = Perm_regdelays_5_3; // @[FFTDesigns.scala 5144:44]
  assign TwiddleFactorsStreamed_clock = clock;
  assign TwiddleFactorsStreamed_reset = reset;
  assign TwiddleFactorsStreamed_io_in_0_Re = PermutationsWithStreaming_1_io_out_0_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_0_Im = PermutationsWithStreaming_1_io_out_0_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_1_Re = PermutationsWithStreaming_1_io_out_1_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_1_Im = PermutationsWithStreaming_1_io_out_1_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_2_Re = PermutationsWithStreaming_1_io_out_2_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_2_Im = PermutationsWithStreaming_1_io_out_2_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_3_Re = PermutationsWithStreaming_1_io_out_3_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_3_Im = PermutationsWithStreaming_1_io_out_3_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_4_Re = PermutationsWithStreaming_1_io_out_4_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_4_Im = PermutationsWithStreaming_1_io_out_4_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_5_Re = PermutationsWithStreaming_1_io_out_5_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_5_Im = PermutationsWithStreaming_1_io_out_5_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_6_Re = PermutationsWithStreaming_1_io_out_6_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_6_Im = PermutationsWithStreaming_1_io_out_6_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_7_Re = PermutationsWithStreaming_1_io_out_7_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_7_Im = PermutationsWithStreaming_1_io_out_7_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_8_Re = PermutationsWithStreaming_1_io_out_8_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_8_Im = PermutationsWithStreaming_1_io_out_8_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_9_Re = PermutationsWithStreaming_1_io_out_9_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_9_Im = PermutationsWithStreaming_1_io_out_9_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_10_Re = PermutationsWithStreaming_1_io_out_10_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_10_Im = PermutationsWithStreaming_1_io_out_10_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_11_Re = PermutationsWithStreaming_1_io_out_11_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_11_Im = PermutationsWithStreaming_1_io_out_11_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_12_Re = PermutationsWithStreaming_1_io_out_12_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_12_Im = PermutationsWithStreaming_1_io_out_12_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_13_Re = PermutationsWithStreaming_1_io_out_13_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_13_Im = PermutationsWithStreaming_1_io_out_13_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_14_Re = PermutationsWithStreaming_1_io_out_14_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_14_Im = PermutationsWithStreaming_1_io_out_14_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_15_Re = PermutationsWithStreaming_1_io_out_15_Re; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_15_Im = PermutationsWithStreaming_1_io_out_15_Im; // @[FFTDesigns.scala 5178:32]
  assign TwiddleFactorsStreamed_io_in_en_0 = Perm_regdelays_1_3; // @[FFTDesigns.scala 5177:38]
  assign TwiddleFactorsStreamed_io_in_en_1 = Twid_regdelays_0_0; // @[FFTDesigns.scala 5186:36]
  assign TwiddleFactorsStreamed_1_clock = clock;
  assign TwiddleFactorsStreamed_1_reset = reset;
  assign TwiddleFactorsStreamed_1_io_in_0_Re = PermutationsWithStreaming_2_io_out_0_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_0_Im = PermutationsWithStreaming_2_io_out_0_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_1_Re = PermutationsWithStreaming_2_io_out_1_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_1_Im = PermutationsWithStreaming_2_io_out_1_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_2_Re = PermutationsWithStreaming_2_io_out_2_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_2_Im = PermutationsWithStreaming_2_io_out_2_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_3_Re = PermutationsWithStreaming_2_io_out_3_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_3_Im = PermutationsWithStreaming_2_io_out_3_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_4_Re = PermutationsWithStreaming_2_io_out_4_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_4_Im = PermutationsWithStreaming_2_io_out_4_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_5_Re = PermutationsWithStreaming_2_io_out_5_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_5_Im = PermutationsWithStreaming_2_io_out_5_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_6_Re = PermutationsWithStreaming_2_io_out_6_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_6_Im = PermutationsWithStreaming_2_io_out_6_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_7_Re = PermutationsWithStreaming_2_io_out_7_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_7_Im = PermutationsWithStreaming_2_io_out_7_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_8_Re = PermutationsWithStreaming_2_io_out_8_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_8_Im = PermutationsWithStreaming_2_io_out_8_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_9_Re = PermutationsWithStreaming_2_io_out_9_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_9_Im = PermutationsWithStreaming_2_io_out_9_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_10_Re = PermutationsWithStreaming_2_io_out_10_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_10_Im = PermutationsWithStreaming_2_io_out_10_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_11_Re = PermutationsWithStreaming_2_io_out_11_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_11_Im = PermutationsWithStreaming_2_io_out_11_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_12_Re = PermutationsWithStreaming_2_io_out_12_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_12_Im = PermutationsWithStreaming_2_io_out_12_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_13_Re = PermutationsWithStreaming_2_io_out_13_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_13_Im = PermutationsWithStreaming_2_io_out_13_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_14_Re = PermutationsWithStreaming_2_io_out_14_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_14_Im = PermutationsWithStreaming_2_io_out_14_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_15_Re = PermutationsWithStreaming_2_io_out_15_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_15_Im = PermutationsWithStreaming_2_io_out_15_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_1_io_in_en_0 = Perm_regdelays_2_3; // @[FFTDesigns.scala 5181:38]
  assign TwiddleFactorsStreamed_1_io_in_en_1 = Twid_regdelays_1_0; // @[FFTDesigns.scala 5186:36]
  assign TwiddleFactorsStreamed_2_clock = clock;
  assign TwiddleFactorsStreamed_2_reset = reset;
  assign TwiddleFactorsStreamed_2_io_in_0_Re = PermutationsWithStreaming_3_io_out_0_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_0_Im = PermutationsWithStreaming_3_io_out_0_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_1_Re = PermutationsWithStreaming_3_io_out_1_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_1_Im = PermutationsWithStreaming_3_io_out_1_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_2_Re = PermutationsWithStreaming_3_io_out_2_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_2_Im = PermutationsWithStreaming_3_io_out_2_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_3_Re = PermutationsWithStreaming_3_io_out_3_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_3_Im = PermutationsWithStreaming_3_io_out_3_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_4_Re = PermutationsWithStreaming_3_io_out_4_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_4_Im = PermutationsWithStreaming_3_io_out_4_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_5_Re = PermutationsWithStreaming_3_io_out_5_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_5_Im = PermutationsWithStreaming_3_io_out_5_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_6_Re = PermutationsWithStreaming_3_io_out_6_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_6_Im = PermutationsWithStreaming_3_io_out_6_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_7_Re = PermutationsWithStreaming_3_io_out_7_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_7_Im = PermutationsWithStreaming_3_io_out_7_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_8_Re = PermutationsWithStreaming_3_io_out_8_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_8_Im = PermutationsWithStreaming_3_io_out_8_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_9_Re = PermutationsWithStreaming_3_io_out_9_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_9_Im = PermutationsWithStreaming_3_io_out_9_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_10_Re = PermutationsWithStreaming_3_io_out_10_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_10_Im = PermutationsWithStreaming_3_io_out_10_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_11_Re = PermutationsWithStreaming_3_io_out_11_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_11_Im = PermutationsWithStreaming_3_io_out_11_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_12_Re = PermutationsWithStreaming_3_io_out_12_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_12_Im = PermutationsWithStreaming_3_io_out_12_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_13_Re = PermutationsWithStreaming_3_io_out_13_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_13_Im = PermutationsWithStreaming_3_io_out_13_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_14_Re = PermutationsWithStreaming_3_io_out_14_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_14_Im = PermutationsWithStreaming_3_io_out_14_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_15_Re = PermutationsWithStreaming_3_io_out_15_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_15_Im = PermutationsWithStreaming_3_io_out_15_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_2_io_in_en_0 = Perm_regdelays_3_3; // @[FFTDesigns.scala 5181:38]
  assign TwiddleFactorsStreamed_2_io_in_en_1 = Twid_regdelays_2_0; // @[FFTDesigns.scala 5186:36]
  assign TwiddleFactorsStreamed_3_clock = clock;
  assign TwiddleFactorsStreamed_3_reset = reset;
  assign TwiddleFactorsStreamed_3_io_in_0_Re = PermutationsWithStreaming_4_io_out_0_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_0_Im = PermutationsWithStreaming_4_io_out_0_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_1_Re = PermutationsWithStreaming_4_io_out_1_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_1_Im = PermutationsWithStreaming_4_io_out_1_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_2_Re = PermutationsWithStreaming_4_io_out_2_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_2_Im = PermutationsWithStreaming_4_io_out_2_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_3_Re = PermutationsWithStreaming_4_io_out_3_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_3_Im = PermutationsWithStreaming_4_io_out_3_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_4_Re = PermutationsWithStreaming_4_io_out_4_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_4_Im = PermutationsWithStreaming_4_io_out_4_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_5_Re = PermutationsWithStreaming_4_io_out_5_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_5_Im = PermutationsWithStreaming_4_io_out_5_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_6_Re = PermutationsWithStreaming_4_io_out_6_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_6_Im = PermutationsWithStreaming_4_io_out_6_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_7_Re = PermutationsWithStreaming_4_io_out_7_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_7_Im = PermutationsWithStreaming_4_io_out_7_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_8_Re = PermutationsWithStreaming_4_io_out_8_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_8_Im = PermutationsWithStreaming_4_io_out_8_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_9_Re = PermutationsWithStreaming_4_io_out_9_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_9_Im = PermutationsWithStreaming_4_io_out_9_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_10_Re = PermutationsWithStreaming_4_io_out_10_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_10_Im = PermutationsWithStreaming_4_io_out_10_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_11_Re = PermutationsWithStreaming_4_io_out_11_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_11_Im = PermutationsWithStreaming_4_io_out_11_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_12_Re = PermutationsWithStreaming_4_io_out_12_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_12_Im = PermutationsWithStreaming_4_io_out_12_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_13_Re = PermutationsWithStreaming_4_io_out_13_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_13_Im = PermutationsWithStreaming_4_io_out_13_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_14_Re = PermutationsWithStreaming_4_io_out_14_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_14_Im = PermutationsWithStreaming_4_io_out_14_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_15_Re = PermutationsWithStreaming_4_io_out_15_Re; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_15_Im = PermutationsWithStreaming_4_io_out_15_Im; // @[FFTDesigns.scala 5182:32]
  assign TwiddleFactorsStreamed_3_io_in_en_0 = Perm_regdelays_4_3; // @[FFTDesigns.scala 5181:38]
  assign TwiddleFactorsStreamed_3_io_in_en_1 = Twid_regdelays_3_0; // @[FFTDesigns.scala 5186:36]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_0_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_0_0 <= Perm_regdelays_0_3; // @[FFTDesigns.scala 5153:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_1_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_1_0 <= Twid_regdelays_0_1; // @[FFTDesigns.scala 5160:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_2_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_2_0 <= Twid_regdelays_1_1; // @[FFTDesigns.scala 5160:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_3_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_3_0 <= Twid_regdelays_2_1; // @[FFTDesigns.scala 5160:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5094:32]
      DFT_regdelays_4_0 <= 1'h0; // @[FFTDesigns.scala 5094:32]
    end else begin
      DFT_regdelays_4_0 <= Twid_regdelays_3_1; // @[FFTDesigns.scala 5160:33]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_0_0 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_0_0 <= Perm_regdelays_1_3; // @[FFTDesigns.scala 5176:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_0_1 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_0_1 <= Twid_regdelays_0_0; // @[FFTDesigns.scala 5185:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_1_0 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_1_0 <= Perm_regdelays_2_3; // @[FFTDesigns.scala 5180:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_1_1 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_1_1 <= Twid_regdelays_1_0; // @[FFTDesigns.scala 5185:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_2_0 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_2_0 <= Perm_regdelays_3_3; // @[FFTDesigns.scala 5180:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_2_1 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_2_1 <= Twid_regdelays_2_0; // @[FFTDesigns.scala 5185:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_3_0 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_3_0 <= Perm_regdelays_4_3; // @[FFTDesigns.scala 5180:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5095:33]
      Twid_regdelays_3_1 <= 1'h0; // @[FFTDesigns.scala 5095:33]
    end else begin
      Twid_regdelays_3_1 <= Twid_regdelays_3_0; // @[FFTDesigns.scala 5185:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_0 <= io_in_ready; // @[FFTDesigns.scala 5122:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_1 <= Perm_regdelays_0_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_2 <= Perm_regdelays_0_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_0_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_0_3 <= Perm_regdelays_0_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_0 <= DFT_regdelays_0_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_1 <= Perm_regdelays_1_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_2 <= Perm_regdelays_1_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_1_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_1_3 <= Perm_regdelays_1_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_0 <= DFT_regdelays_1_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_1 <= Perm_regdelays_2_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_2 <= Perm_regdelays_2_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_2_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_2_3 <= Perm_regdelays_2_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_0 <= DFT_regdelays_2_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_1 <= Perm_regdelays_3_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_2 <= Perm_regdelays_3_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_3_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_3_3 <= Perm_regdelays_3_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_0 <= DFT_regdelays_3_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_1 <= Perm_regdelays_4_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_2 <= Perm_regdelays_4_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_4_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_4_3 <= Perm_regdelays_4_2; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_0 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_0 <= DFT_regdelays_4_0; // @[FFTDesigns.scala 5132:34]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_1 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_1 <= Perm_regdelays_5_0; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_2 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_2 <= Perm_regdelays_5_1; // @[FFTDesigns.scala 5141:32]
    end
    if (reset) begin // @[FFTDesigns.scala 5096:33]
      Perm_regdelays_5_3 <= 1'h0; // @[FFTDesigns.scala 5096:33]
    end else begin
      Perm_regdelays_5_3 <= Perm_regdelays_5_2; // @[FFTDesigns.scala 5141:32]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DFT_regdelays_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  DFT_regdelays_1_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  DFT_regdelays_2_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  DFT_regdelays_3_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  DFT_regdelays_4_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  Twid_regdelays_0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  Twid_regdelays_0_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  Twid_regdelays_1_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  Twid_regdelays_1_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  Twid_regdelays_2_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  Twid_regdelays_2_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  Twid_regdelays_3_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  Twid_regdelays_3_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  Perm_regdelays_0_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  Perm_regdelays_0_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  Perm_regdelays_0_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  Perm_regdelays_0_3 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  Perm_regdelays_1_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  Perm_regdelays_1_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  Perm_regdelays_1_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  Perm_regdelays_1_3 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  Perm_regdelays_2_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  Perm_regdelays_2_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  Perm_regdelays_2_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  Perm_regdelays_2_3 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  Perm_regdelays_3_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  Perm_regdelays_3_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  Perm_regdelays_3_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  Perm_regdelays_3_3 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  Perm_regdelays_4_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  Perm_regdelays_4_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  Perm_regdelays_4_2 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  Perm_regdelays_4_3 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  Perm_regdelays_5_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  Perm_regdelays_5_1 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  Perm_regdelays_5_2 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  Perm_regdelays_5_3 = _RAND_36[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexSub(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  input  [31:0] io_in_b_Re,
  input  [31:0] io_in_b_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire  FP_subber_clock; // @[FPComplex.scala 78:25]
  wire  FP_subber_reset; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_in_a; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_in_b; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_io_out_s; // @[FPComplex.scala 78:25]
  wire  FP_subber_1_clock; // @[FPComplex.scala 78:25]
  wire  FP_subber_1_reset; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_in_a; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_in_b; // @[FPComplex.scala 78:25]
  wire [31:0] FP_subber_1_io_out_s; // @[FPComplex.scala 78:25]
  FP_subber FP_subber ( // @[FPComplex.scala 78:25]
    .clock(FP_subber_clock),
    .reset(FP_subber_reset),
    .io_in_a(FP_subber_io_in_a),
    .io_in_b(FP_subber_io_in_b),
    .io_out_s(FP_subber_io_out_s)
  );
  FP_subber FP_subber_1 ( // @[FPComplex.scala 78:25]
    .clock(FP_subber_1_clock),
    .reset(FP_subber_1_reset),
    .io_in_a(FP_subber_1_io_in_a),
    .io_in_b(FP_subber_1_io_in_b),
    .io_out_s(FP_subber_1_io_out_s)
  );
  assign io_out_s_Re = FP_subber_io_out_s; // @[FPComplex.scala 85:17]
  assign io_out_s_Im = FP_subber_1_io_out_s; // @[FPComplex.scala 86:17]
  assign FP_subber_clock = clock;
  assign FP_subber_reset = reset;
  assign FP_subber_io_in_a = io_in_a_Re; // @[FPComplex.scala 81:24]
  assign FP_subber_io_in_b = io_in_b_Re; // @[FPComplex.scala 82:24]
  assign FP_subber_1_clock = clock;
  assign FP_subber_1_reset = reset;
  assign FP_subber_1_io_in_a = io_in_a_Im; // @[FPComplex.scala 83:24]
  assign FP_subber_1_io_in_b = io_in_b_Im; // @[FPComplex.scala 84:24]
endmodule
module FPComplexMultiAdder_80(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  output [31:0] io_out_Re,
  output [31:0] io_out_Im
);
  assign io_out_Re = io_in_0_Re; // @[FPComplex.scala 521:14]
  assign io_out_Im = io_in_0_Im; // @[FPComplex.scala 521:14]
endmodule
module FPComplexMult_reducable_v2(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 380:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 380:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 380:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 380:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 380:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 380:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 380:33]
  reg [31:0] result_0_Re; // @[FPComplex.scala 391:31]
  reg [31:0] result_0_Im; // @[FPComplex.scala 391:31]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 380:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  assign io_out_s_Re = result_0_Re; // @[FPComplex.scala 400:20]
  assign io_out_s_Im = result_0_Im; // @[FPComplex.scala 400:20]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 381:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 381:24]
  assign cmplx_adj_io_in_adj = 8'h1; // @[FPComplex.scala 384:30]
  assign cmplx_adj_io_is_neg = 1'h1; // @[FPComplex.scala 386:32]
  assign cmplx_adj_io_is_flip = 1'h0; // @[FPComplex.scala 382:29]
  always @(posedge clock) begin
    if (reset) begin // @[FPComplex.scala 391:31]
      result_0_Re <= 32'h0; // @[FPComplex.scala 391:31]
    end else begin
      result_0_Re <= cmplx_adj_io_out_Re; // @[FPComplex.scala 394:25]
    end
    if (reset) begin // @[FPComplex.scala 391:31]
      result_0_Im <= 32'h0; // @[FPComplex.scala 391:31]
    end else begin
      result_0_Im <= cmplx_adj_io_out_Im; // @[FPComplex.scala 394:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  result_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  result_0_Im = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FPComplexMult_reducable_v2_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_Re,
  input  [31:0] io_in_a_Im,
  output [31:0] io_out_s_Re,
  output [31:0] io_out_s_Im
);
  wire [31:0] cmplx_adj_io_in_Re; // @[FPComplex.scala 340:33]
  wire [31:0] cmplx_adj_io_in_Im; // @[FPComplex.scala 340:33]
  wire [7:0] cmplx_adj_io_in_adj; // @[FPComplex.scala 340:33]
  wire  cmplx_adj_io_is_neg; // @[FPComplex.scala 340:33]
  wire  cmplx_adj_io_is_flip; // @[FPComplex.scala 340:33]
  wire [31:0] cmplx_adj_io_out_Re; // @[FPComplex.scala 340:33]
  wire [31:0] cmplx_adj_io_out_Im; // @[FPComplex.scala 340:33]
  wire  FP_multiplier_clock; // @[FPComplex.scala 368:29]
  wire  FP_multiplier_reset; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_io_in_a; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_io_in_b; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_io_out_s; // @[FPComplex.scala 368:29]
  wire  FP_multiplier_1_clock; // @[FPComplex.scala 368:29]
  wire  FP_multiplier_1_reset; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_1_io_in_a; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_1_io_in_b; // @[FPComplex.scala 368:29]
  wire [31:0] FP_multiplier_1_io_out_s; // @[FPComplex.scala 368:29]
  cmplx_adj cmplx_adj ( // @[FPComplex.scala 340:33]
    .io_in_Re(cmplx_adj_io_in_Re),
    .io_in_Im(cmplx_adj_io_in_Im),
    .io_in_adj(cmplx_adj_io_in_adj),
    .io_is_neg(cmplx_adj_io_is_neg),
    .io_is_flip(cmplx_adj_io_is_flip),
    .io_out_Re(cmplx_adj_io_out_Re),
    .io_out_Im(cmplx_adj_io_out_Im)
  );
  FP_multiplier FP_multiplier ( // @[FPComplex.scala 368:29]
    .clock(FP_multiplier_clock),
    .reset(FP_multiplier_reset),
    .io_in_a(FP_multiplier_io_in_a),
    .io_in_b(FP_multiplier_io_in_b),
    .io_out_s(FP_multiplier_io_out_s)
  );
  FP_multiplier FP_multiplier_1 ( // @[FPComplex.scala 368:29]
    .clock(FP_multiplier_1_clock),
    .reset(FP_multiplier_1_reset),
    .io_in_a(FP_multiplier_1_io_in_a),
    .io_in_b(FP_multiplier_1_io_in_b),
    .io_out_s(FP_multiplier_1_io_out_s)
  );
  assign io_out_s_Re = FP_multiplier_io_out_s; // @[FPComplex.scala 375:21]
  assign io_out_s_Im = FP_multiplier_1_io_out_s; // @[FPComplex.scala 376:21]
  assign cmplx_adj_io_in_Re = io_in_a_Re; // @[FPComplex.scala 341:24]
  assign cmplx_adj_io_in_Im = io_in_a_Im; // @[FPComplex.scala 341:24]
  assign cmplx_adj_io_in_adj = 8'h0; // @[FPComplex.scala 365:30]
  assign cmplx_adj_io_is_neg = 1'h0; // @[FPComplex.scala 366:30]
  assign cmplx_adj_io_is_flip = 1'h1; // @[FPComplex.scala 342:29]
  assign FP_multiplier_clock = clock;
  assign FP_multiplier_reset = reset;
  assign FP_multiplier_io_in_a = cmplx_adj_io_out_Re; // @[FPComplex.scala 371:29]
  assign FP_multiplier_io_in_b = 32'hbf5db3d6; // @[FPComplex.scala 372:29]
  assign FP_multiplier_1_clock = clock;
  assign FP_multiplier_1_reset = reset;
  assign FP_multiplier_1_io_in_a = cmplx_adj_io_out_Im; // @[FPComplex.scala 373:29]
  assign FP_multiplier_1_io_in_b = 32'hbf5db3d6; // @[FPComplex.scala 374:29]
endmodule
module DFT_r_v2_40(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  FPComplexAdder_clock; // @[FFTDesigns.scala 258:34]
  wire  FPComplexAdder_reset; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_a_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_a_Im; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_b_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_in_b_Im; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 258:34]
  wire [31:0] FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 258:34]
  wire  FPComplexSub_clock; // @[FFTDesigns.scala 261:34]
  wire  FPComplexSub_reset; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_a_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_a_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_b_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_in_b_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_out_s_Re; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexSub_io_out_s_Im; // @[FFTDesigns.scala 261:34]
  wire [31:0] FPComplexMultiAdder_io_in_0_Re; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_in_0_Im; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 275:36]
  wire [31:0] FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 275:36]
  wire  FPComplexMult_reducable_v2_clock; // @[FFTDesigns.scala 294:39]
  wire  FPComplexMult_reducable_v2_reset; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Re; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_in_a_Im; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 294:39]
  wire [31:0] FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 294:39]
  wire  FPComplexMult_reducable_v2_1_clock; // @[FFTDesigns.scala 297:39]
  wire  FPComplexMult_reducable_v2_1_reset; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Re; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_in_a_Im; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 297:39]
  wire [31:0] FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 297:39]
  wire  FPComplexAdder_reducable_clock; // @[FFTDesigns.scala 338:34]
  wire  FPComplexAdder_reducable_reset; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_a_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_a_Im; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_b_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_in_b_Im; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_out_s_Re; // @[FFTDesigns.scala 338:34]
  wire [31:0] FPComplexAdder_reducable_io_out_s_Im; // @[FFTDesigns.scala 338:34]
  wire  FPComplexSub_reducable_clock; // @[FFTDesigns.scala 341:34]
  wire  FPComplexSub_reducable_reset; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_a_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_a_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_b_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_in_b_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_out_s_Re; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexSub_reducable_io_out_s_Im; // @[FFTDesigns.scala 341:34]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_in_0_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_in_0_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_in_0_Im; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_out_Re; // @[FFTDesigns.scala 394:29]
  wire [31:0] FPComplexMultiAdder_2_io_out_Im; // @[FFTDesigns.scala 394:29]
  wire  FPComplexAdder_1_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_1_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_1_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_2_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_2_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_2_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_3_clock; // @[FFTDesigns.scala 418:27]
  wire  FPComplexAdder_3_reset; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_a_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_a_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_b_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_in_b_Im; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_out_s_Re; // @[FFTDesigns.scala 418:27]
  wire [31:0] FPComplexAdder_3_io_out_s_Im; // @[FFTDesigns.scala 418:27]
  reg [31:0] initial_layer_out_0_0_Re; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_0_0_Im; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_1_0_Re; // @[FFTDesigns.scala 276:84]
  reg [31:0] initial_layer_out_1_0_Im; // @[FFTDesigns.scala 276:84]
  reg [31:0] finallayer_0_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_0_Im; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_1_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_1_Im; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_2_Re; // @[FFTDesigns.scala 421:31]
  reg [31:0] finallayer_2_Im; // @[FFTDesigns.scala 421:31]
  FPComplexAdder FPComplexAdder ( // @[FFTDesigns.scala 258:34]
    .clock(FPComplexAdder_clock),
    .reset(FPComplexAdder_reset),
    .io_in_a_Re(FPComplexAdder_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_io_out_s_Im)
  );
  FPComplexSub FPComplexSub ( // @[FFTDesigns.scala 261:34]
    .clock(FPComplexSub_clock),
    .reset(FPComplexSub_reset),
    .io_in_a_Re(FPComplexSub_io_in_a_Re),
    .io_in_a_Im(FPComplexSub_io_in_a_Im),
    .io_in_b_Re(FPComplexSub_io_in_b_Re),
    .io_in_b_Im(FPComplexSub_io_in_b_Im),
    .io_out_s_Re(FPComplexSub_io_out_s_Re),
    .io_out_s_Im(FPComplexSub_io_out_s_Im)
  );
  FPComplexMultiAdder_80 FPComplexMultiAdder ( // @[FFTDesigns.scala 275:36]
    .io_in_0_Re(FPComplexMultiAdder_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_io_out_Im)
  );
  FPComplexMult_reducable_v2 FPComplexMult_reducable_v2 ( // @[FFTDesigns.scala 294:39]
    .clock(FPComplexMult_reducable_v2_clock),
    .reset(FPComplexMult_reducable_v2_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_io_out_s_Im)
  );
  FPComplexMult_reducable_v2_1 FPComplexMult_reducable_v2_1 ( // @[FFTDesigns.scala 297:39]
    .clock(FPComplexMult_reducable_v2_1_clock),
    .reset(FPComplexMult_reducable_v2_1_reset),
    .io_in_a_Re(FPComplexMult_reducable_v2_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_reducable_v2_1_io_in_a_Im),
    .io_out_s_Re(FPComplexMult_reducable_v2_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_reducable_v2_1_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_reducable ( // @[FFTDesigns.scala 338:34]
    .clock(FPComplexAdder_reducable_clock),
    .reset(FPComplexAdder_reducable_reset),
    .io_in_a_Re(FPComplexAdder_reducable_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_reducable_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_reducable_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_reducable_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_reducable_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_reducable_io_out_s_Im)
  );
  FPComplexSub FPComplexSub_reducable ( // @[FFTDesigns.scala 341:34]
    .clock(FPComplexSub_reducable_clock),
    .reset(FPComplexSub_reducable_reset),
    .io_in_a_Re(FPComplexSub_reducable_io_in_a_Re),
    .io_in_a_Im(FPComplexSub_reducable_io_in_a_Im),
    .io_in_b_Re(FPComplexSub_reducable_io_in_b_Re),
    .io_in_b_Im(FPComplexSub_reducable_io_in_b_Im),
    .io_out_s_Re(FPComplexSub_reducable_io_out_s_Re),
    .io_out_s_Im(FPComplexSub_reducable_io_out_s_Im)
  );
  FPComplexMultiAdder_80 FPComplexMultiAdder_1 ( // @[FFTDesigns.scala 394:29]
    .io_in_0_Re(FPComplexMultiAdder_1_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_1_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_1_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_1_io_out_Im)
  );
  FPComplexMultiAdder_80 FPComplexMultiAdder_2 ( // @[FFTDesigns.scala 394:29]
    .io_in_0_Re(FPComplexMultiAdder_2_io_in_0_Re),
    .io_in_0_Im(FPComplexMultiAdder_2_io_in_0_Im),
    .io_out_Re(FPComplexMultiAdder_2_io_out_Re),
    .io_out_Im(FPComplexMultiAdder_2_io_out_Im)
  );
  FPComplexAdder FPComplexAdder_1 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_1_clock),
    .reset(FPComplexAdder_1_reset),
    .io_in_a_Re(FPComplexAdder_1_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_1_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_1_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_1_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_1_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_1_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_2 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_2_clock),
    .reset(FPComplexAdder_2_reset),
    .io_in_a_Re(FPComplexAdder_2_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_2_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_2_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_2_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_2_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_2_io_out_s_Im)
  );
  FPComplexAdder FPComplexAdder_3 ( // @[FFTDesigns.scala 418:27]
    .clock(FPComplexAdder_3_clock),
    .reset(FPComplexAdder_3_reset),
    .io_in_a_Re(FPComplexAdder_3_io_in_a_Re),
    .io_in_a_Im(FPComplexAdder_3_io_in_a_Im),
    .io_in_b_Re(FPComplexAdder_3_io_in_b_Re),
    .io_in_b_Im(FPComplexAdder_3_io_in_b_Im),
    .io_out_s_Re(FPComplexAdder_3_io_out_s_Re),
    .io_out_s_Im(FPComplexAdder_3_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexAdder_1_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_0_Im = FPComplexAdder_1_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign io_out_1_Re = FPComplexAdder_2_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_1_Im = FPComplexAdder_2_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign io_out_2_Re = FPComplexAdder_3_io_out_s_Re; // @[FFTDesigns.scala 432:19]
  assign io_out_2_Im = FPComplexAdder_3_io_out_s_Im; // @[FFTDesigns.scala 432:19]
  assign FPComplexAdder_clock = clock;
  assign FPComplexAdder_reset = reset;
  assign FPComplexAdder_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 268:38]
  assign FPComplexAdder_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 268:38]
  assign FPComplexAdder_io_in_b_Re = io_in_2_Re; // @[FFTDesigns.scala 269:38]
  assign FPComplexAdder_io_in_b_Im = io_in_2_Im; // @[FFTDesigns.scala 269:38]
  assign FPComplexSub_clock = clock;
  assign FPComplexSub_reset = reset;
  assign FPComplexSub_io_in_a_Re = io_in_1_Re; // @[FFTDesigns.scala 270:38]
  assign FPComplexSub_io_in_a_Im = io_in_1_Im; // @[FFTDesigns.scala 270:38]
  assign FPComplexSub_io_in_b_Re = io_in_2_Re; // @[FFTDesigns.scala 271:38]
  assign FPComplexSub_io_in_b_Im = io_in_2_Im; // @[FFTDesigns.scala 271:38]
  assign FPComplexMultiAdder_io_in_0_Re = initial_layer_out_1_0_Re; // @[FFTDesigns.scala 290:27]
  assign FPComplexMultiAdder_io_in_0_Im = initial_layer_out_1_0_Im; // @[FFTDesigns.scala 290:27]
  assign FPComplexMult_reducable_v2_clock = clock;
  assign FPComplexMult_reducable_v2_reset = reset;
  assign FPComplexMult_reducable_v2_io_in_a_Re = FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 320:34]
  assign FPComplexMult_reducable_v2_io_in_a_Im = FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 320:34]
  assign FPComplexMult_reducable_v2_1_clock = clock;
  assign FPComplexMult_reducable_v2_1_reset = reset;
  assign FPComplexMult_reducable_v2_1_io_in_a_Re = FPComplexSub_io_out_s_Re; // @[FFTDesigns.scala 323:34]
  assign FPComplexMult_reducable_v2_1_io_in_a_Im = FPComplexSub_io_out_s_Im; // @[FFTDesigns.scala 323:34]
  assign FPComplexAdder_reducable_clock = clock;
  assign FPComplexAdder_reducable_reset = reset;
  assign FPComplexAdder_reducable_io_in_a_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 366:36]
  assign FPComplexAdder_reducable_io_in_a_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 366:36]
  assign FPComplexAdder_reducable_io_in_b_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 367:36]
  assign FPComplexAdder_reducable_io_in_b_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 367:36]
  assign FPComplexSub_reducable_clock = clock;
  assign FPComplexSub_reducable_reset = reset;
  assign FPComplexSub_reducable_io_in_a_Re = FPComplexMult_reducable_v2_io_out_s_Re; // @[FFTDesigns.scala 368:36]
  assign FPComplexSub_reducable_io_in_a_Im = FPComplexMult_reducable_v2_io_out_s_Im; // @[FFTDesigns.scala 368:36]
  assign FPComplexSub_reducable_io_in_b_Re = FPComplexMult_reducable_v2_1_io_out_s_Re; // @[FFTDesigns.scala 369:36]
  assign FPComplexSub_reducable_io_in_b_Im = FPComplexMult_reducable_v2_1_io_out_s_Im; // @[FFTDesigns.scala 369:36]
  assign FPComplexMultiAdder_1_io_in_0_Re = FPComplexAdder_reducable_io_out_s_Re; // @[FFTDesigns.scala 402:36]
  assign FPComplexMultiAdder_1_io_in_0_Im = FPComplexAdder_reducable_io_out_s_Im; // @[FFTDesigns.scala 402:36]
  assign FPComplexMultiAdder_2_io_in_0_Re = FPComplexSub_reducable_io_out_s_Re; // @[FFTDesigns.scala 404:61]
  assign FPComplexMultiAdder_2_io_in_0_Im = FPComplexSub_reducable_io_out_s_Im; // @[FFTDesigns.scala 404:61]
  assign FPComplexAdder_1_clock = clock;
  assign FPComplexAdder_1_reset = reset;
  assign FPComplexAdder_1_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_1_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_1_io_in_b_Re = FPComplexMultiAdder_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_1_io_in_b_Im = FPComplexMultiAdder_io_out_Im; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_2_clock = clock;
  assign FPComplexAdder_2_reset = reset;
  assign FPComplexAdder_2_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_2_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_2_io_in_b_Re = FPComplexMultiAdder_1_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_2_io_in_b_Im = FPComplexMultiAdder_1_io_out_Im; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_3_clock = clock;
  assign FPComplexAdder_3_reset = reset;
  assign FPComplexAdder_3_io_in_a_Re = finallayer_2_Re; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_3_io_in_a_Im = finallayer_2_Im; // @[FFTDesigns.scala 430:35]
  assign FPComplexAdder_3_io_in_b_Re = FPComplexMultiAdder_2_io_out_Re; // @[FFTDesigns.scala 431:35]
  assign FPComplexAdder_3_io_in_b_Im = FPComplexMultiAdder_2_io_out_Im; // @[FFTDesigns.scala 431:35]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_0_0_Re <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_0_0_Re <= FPComplexAdder_io_out_s_Re; // @[FFTDesigns.scala 281:37]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_0_0_Im <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_0_0_Im <= FPComplexAdder_io_out_s_Im; // @[FFTDesigns.scala 281:37]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_1_0_Re <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_1_0_Re <= initial_layer_out_0_0_Re; // @[FFTDesigns.scala 284:32]
    end
    if (reset) begin // @[FFTDesigns.scala 276:84]
      initial_layer_out_1_0_Im <= 32'h0; // @[FFTDesigns.scala 276:84]
    end else begin
      initial_layer_out_1_0_Im <= initial_layer_out_0_0_Im; // @[FFTDesigns.scala 284:32]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_0_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_0_Re <= io_in_0_Re; // @[FFTDesigns.scala 424:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_0_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_0_Im <= io_in_0_Im; // @[FFTDesigns.scala 424:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_1_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_1_Re <= finallayer_0_Re; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_1_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_1_Im <= finallayer_0_Im; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_2_Re <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_2_Re <= finallayer_1_Re; // @[FFTDesigns.scala 426:25]
    end
    if (reset) begin // @[FFTDesigns.scala 421:31]
      finallayer_2_Im <= 32'h0; // @[FFTDesigns.scala 421:31]
    end else begin
      finallayer_2_Im <= finallayer_1_Im; // @[FFTDesigns.scala 426:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  initial_layer_out_0_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  initial_layer_out_0_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  initial_layer_out_1_0_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  initial_layer_out_1_0_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  finallayer_0_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  finallayer_0_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  finallayer_1_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  finallayer_1_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  finallayer_2_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  finallayer_2_Im = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_Block_192(
  input         clock,
  input  [3:0]  io_in_raddr,
  input  [3:0]  io_in_waddr,
  input  [31:0] io_in_data_Re,
  input  [31:0] io_in_data_Im,
  input         io_re,
  input         io_wr,
  input         io_en,
  output [31:0] io_out_data_Re,
  output [31:0] io_out_data_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_0_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_8_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_8_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_9_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_9_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_10_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_10_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_11_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_11_Im; // @[FFTDesigns.scala 3286:18]
  wire [31:0] _GEN_49 = 4'h1 == io_in_raddr ? mem_1_Im : mem_0_Im; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_50 = 4'h2 == io_in_raddr ? mem_2_Im : _GEN_49; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_51 = 4'h3 == io_in_raddr ? mem_3_Im : _GEN_50; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_52 = 4'h4 == io_in_raddr ? mem_4_Im : _GEN_51; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_53 = 4'h5 == io_in_raddr ? mem_5_Im : _GEN_52; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_54 = 4'h6 == io_in_raddr ? mem_6_Im : _GEN_53; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_55 = 4'h7 == io_in_raddr ? mem_7_Im : _GEN_54; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_56 = 4'h8 == io_in_raddr ? mem_8_Im : _GEN_55; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_57 = 4'h9 == io_in_raddr ? mem_9_Im : _GEN_56; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_58 = 4'ha == io_in_raddr ? mem_10_Im : _GEN_57; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_59 = 4'hb == io_in_raddr ? mem_11_Im : _GEN_58; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_61 = 4'h1 == io_in_raddr ? mem_1_Re : mem_0_Re; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_62 = 4'h2 == io_in_raddr ? mem_2_Re : _GEN_61; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_63 = 4'h3 == io_in_raddr ? mem_3_Re : _GEN_62; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_64 = 4'h4 == io_in_raddr ? mem_4_Re : _GEN_63; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_65 = 4'h5 == io_in_raddr ? mem_5_Re : _GEN_64; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_66 = 4'h6 == io_in_raddr ? mem_6_Re : _GEN_65; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_67 = 4'h7 == io_in_raddr ? mem_7_Re : _GEN_66; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_68 = 4'h8 == io_in_raddr ? mem_8_Re : _GEN_67; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_69 = 4'h9 == io_in_raddr ? mem_9_Re : _GEN_68; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_70 = 4'ha == io_in_raddr ? mem_10_Re : _GEN_69; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_71 = 4'hb == io_in_raddr ? mem_11_Re : _GEN_70; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_72 = io_re ? _GEN_59 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3295:24]
  wire [31:0] _GEN_73 = io_re ? _GEN_71 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3294:24]
  assign io_out_data_Re = io_en ? _GEN_73 : 32'h0; // @[FFTDesigns.scala 3287:16 3298:22]
  assign io_out_data_Im = io_en ? _GEN_72 : 32'h0; // @[FFTDesigns.scala 3287:16 3299:22]
  always @(posedge clock) begin
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h8 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_8_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h8 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_8_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h9 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_9_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'h9 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_9_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'ha == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_10_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'ha == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_10_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hb == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_11_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (4'hb == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_11_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_3_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_4_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_4_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_5_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_5_Im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_6_Re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_6_Im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_7_Re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_7_Im = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mem_8_Re = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mem_8_Im = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_9_Re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mem_9_Im = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mem_10_Re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mem_10_Im = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_11_Re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mem_11_Im = _RAND_23[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module M0_Config_ROM_6(
  input  [2:0] io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11,
  output [3:0] io_out_12,
  output [3:0] io_out_13,
  output [3:0] io_out_14,
  output [3:0] io_out_15
);
  wire [3:0] _GEN_1 = 3'h1 == io_in_cnt ? 4'h1 : 4'h0; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_2 = 3'h2 == io_in_cnt ? 4'h2 : _GEN_1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_3 = 3'h3 == io_in_cnt ? 4'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_4 = 3'h4 == io_in_cnt ? 4'h4 : _GEN_3; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_7 = 3'h1 == io_in_cnt ? 4'h3 : 4'h2; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_8 = 3'h2 == io_in_cnt ? 4'h4 : _GEN_7; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_9 = 3'h3 == io_in_cnt ? 4'h5 : _GEN_8; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_10 = 3'h4 == io_in_cnt ? 4'h0 : _GEN_9; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_13 = 3'h1 == io_in_cnt ? 4'h2 : 4'h1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_14 = 3'h2 == io_in_cnt ? 4'h3 : _GEN_13; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_15 = 3'h3 == io_in_cnt ? 4'h4 : _GEN_14; // @[FFTDesigns.scala 3227:{17,17}]
  wire [3:0] _GEN_16 = 3'h4 == io_in_cnt ? 4'h5 : _GEN_15; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_0 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_4; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_1 = 3'h5 == io_in_cnt ? 4'h1 : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_2 = 3'h5 == io_in_cnt ? 4'h0 : _GEN_16; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_3 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_4; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_4 = 3'h5 == io_in_cnt ? 4'h1 : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_5 = 3'h5 == io_in_cnt ? 4'h0 : _GEN_16; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_6 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_4; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_7 = 3'h5 == io_in_cnt ? 4'h1 : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_8 = 3'h5 == io_in_cnt ? 4'h0 : _GEN_16; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_9 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_4; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_10 = 3'h5 == io_in_cnt ? 4'h1 : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_11 = 3'h5 == io_in_cnt ? 4'h0 : _GEN_16; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_12 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_4; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_13 = 3'h5 == io_in_cnt ? 4'h1 : _GEN_10; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_14 = 3'h5 == io_in_cnt ? 4'h0 : _GEN_16; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_15 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_4; // @[FFTDesigns.scala 3227:{17,17}]
endmodule
module M1_Config_ROM_6(
  input  [2:0] io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11,
  output [3:0] io_out_12,
  output [3:0] io_out_13,
  output [3:0] io_out_14,
  output [3:0] io_out_15
);
  wire [3:0] _GEN_1 = 3'h1 == io_in_cnt ? 4'h3 : 4'h0; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_2 = 3'h2 == io_in_cnt ? 4'h5 : _GEN_1; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_3 = 3'h3 == io_in_cnt ? 4'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_4 = 3'h4 == io_in_cnt ? 4'h2 : _GEN_3; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_31 = 3'h1 == io_in_cnt ? 4'h2 : 4'h0; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_32 = 3'h2 == io_in_cnt ? 4'h5 : _GEN_31; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_33 = 3'h3 == io_in_cnt ? 4'h1 : _GEN_32; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_34 = 3'h4 == io_in_cnt ? 4'h3 : _GEN_33; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_62 = 3'h2 == io_in_cnt ? 4'h4 : _GEN_31; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_63 = 3'h3 == io_in_cnt ? 4'h1 : _GEN_62; // @[FFTDesigns.scala 3250:{17,17}]
  wire [3:0] _GEN_64 = 3'h4 == io_in_cnt ? 4'h3 : _GEN_63; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_0 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_4; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_1 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_4; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_2 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_4; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_3 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_4; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_4 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_4; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_5 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_34; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_6 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_34; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_7 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_34; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_8 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_34; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_9 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_34; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_10 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_64; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_11 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_64; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_12 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_64; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_13 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_64; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_14 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_64; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_15 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_64; // @[FFTDesigns.scala 3250:{17,17}]
endmodule
module Streaming_Permute_Config_6(
  input  [2:0] io_in_cnt,
  output [3:0] io_out_0,
  output [3:0] io_out_1,
  output [3:0] io_out_2,
  output [3:0] io_out_3,
  output [3:0] io_out_4,
  output [3:0] io_out_5,
  output [3:0] io_out_6,
  output [3:0] io_out_7,
  output [3:0] io_out_8,
  output [3:0] io_out_9,
  output [3:0] io_out_10,
  output [3:0] io_out_11,
  output [3:0] io_out_12,
  output [3:0] io_out_13,
  output [3:0] io_out_14
);
  wire [3:0] _GEN_1 = 3'h1 == io_in_cnt ? 4'h5 : 4'h0; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_2 = 3'h2 == io_in_cnt ? 4'ha : _GEN_1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_3 = 3'h3 == io_in_cnt ? 4'h0 : _GEN_2; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_4 = 3'h4 == io_in_cnt ? 4'h5 : _GEN_3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_7 = 3'h1 == io_in_cnt ? 4'h0 : 4'hb; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_8 = 3'h2 == io_in_cnt ? 4'h5 : _GEN_7; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_9 = 3'h3 == io_in_cnt ? 4'hb : _GEN_8; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_10 = 3'h4 == io_in_cnt ? 4'h0 : _GEN_9; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_13 = 3'h1 == io_in_cnt ? 4'hb : 4'h6; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_14 = 3'h2 == io_in_cnt ? 4'h0 : _GEN_13; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_15 = 3'h3 == io_in_cnt ? 4'h6 : _GEN_14; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_16 = 3'h4 == io_in_cnt ? 4'hb : _GEN_15; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_19 = 3'h1 == io_in_cnt ? 4'h6 : 4'h1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_20 = 3'h2 == io_in_cnt ? 4'hb : _GEN_19; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_21 = 3'h3 == io_in_cnt ? 4'h1 : _GEN_20; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_22 = 3'h4 == io_in_cnt ? 4'h6 : _GEN_21; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_25 = 3'h1 == io_in_cnt ? 4'h1 : 4'hc; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_26 = 3'h2 == io_in_cnt ? 4'h6 : _GEN_25; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_27 = 3'h3 == io_in_cnt ? 4'hc : _GEN_26; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_28 = 3'h4 == io_in_cnt ? 4'h1 : _GEN_27; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_31 = 3'h1 == io_in_cnt ? 4'hc : 4'h7; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_32 = 3'h2 == io_in_cnt ? 4'h1 : _GEN_31; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_33 = 3'h3 == io_in_cnt ? 4'h7 : _GEN_32; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_34 = 3'h4 == io_in_cnt ? 4'hc : _GEN_33; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_37 = 3'h1 == io_in_cnt ? 4'h7 : 4'h2; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_38 = 3'h2 == io_in_cnt ? 4'hc : _GEN_37; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_39 = 3'h3 == io_in_cnt ? 4'h2 : _GEN_38; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_40 = 3'h4 == io_in_cnt ? 4'h7 : _GEN_39; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_43 = 3'h1 == io_in_cnt ? 4'h2 : 4'hd; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_44 = 3'h2 == io_in_cnt ? 4'h7 : _GEN_43; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_45 = 3'h3 == io_in_cnt ? 4'hd : _GEN_44; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_46 = 3'h4 == io_in_cnt ? 4'h2 : _GEN_45; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_49 = 3'h1 == io_in_cnt ? 4'hd : 4'h8; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_50 = 3'h2 == io_in_cnt ? 4'h2 : _GEN_49; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_51 = 3'h3 == io_in_cnt ? 4'h8 : _GEN_50; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_52 = 3'h4 == io_in_cnt ? 4'hd : _GEN_51; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_55 = 3'h1 == io_in_cnt ? 4'h8 : 4'h3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_56 = 3'h2 == io_in_cnt ? 4'hd : _GEN_55; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_57 = 3'h3 == io_in_cnt ? 4'h3 : _GEN_56; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_58 = 3'h4 == io_in_cnt ? 4'h8 : _GEN_57; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_61 = 3'h1 == io_in_cnt ? 4'h3 : 4'he; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_62 = 3'h2 == io_in_cnt ? 4'h8 : _GEN_61; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_63 = 3'h3 == io_in_cnt ? 4'he : _GEN_62; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_64 = 3'h4 == io_in_cnt ? 4'h3 : _GEN_63; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_67 = 3'h1 == io_in_cnt ? 4'he : 4'h9; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_68 = 3'h2 == io_in_cnt ? 4'h3 : _GEN_67; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_69 = 3'h3 == io_in_cnt ? 4'h9 : _GEN_68; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_70 = 3'h4 == io_in_cnt ? 4'he : _GEN_69; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_73 = 3'h1 == io_in_cnt ? 4'h9 : 4'h4; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_74 = 3'h2 == io_in_cnt ? 4'he : _GEN_73; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_75 = 3'h3 == io_in_cnt ? 4'h4 : _GEN_74; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_76 = 3'h4 == io_in_cnt ? 4'h9 : _GEN_75; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_79 = 3'h1 == io_in_cnt ? 4'h4 : 4'hf; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_80 = 3'h2 == io_in_cnt ? 4'h9 : _GEN_79; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_81 = 3'h3 == io_in_cnt ? 4'hf : _GEN_80; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_82 = 3'h4 == io_in_cnt ? 4'h4 : _GEN_81; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_85 = 3'h1 == io_in_cnt ? 4'hf : 4'ha; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_86 = 3'h2 == io_in_cnt ? 4'h4 : _GEN_85; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_87 = 3'h3 == io_in_cnt ? 4'ha : _GEN_86; // @[FFTDesigns.scala 3273:{17,17}]
  wire [3:0] _GEN_88 = 3'h4 == io_in_cnt ? 4'hf : _GEN_87; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_0 = 3'h5 == io_in_cnt ? 4'ha : _GEN_4; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_1 = 3'h5 == io_in_cnt ? 4'h5 : _GEN_10; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_2 = 3'h5 == io_in_cnt ? 4'h0 : _GEN_16; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_3 = 3'h5 == io_in_cnt ? 4'hb : _GEN_22; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_4 = 3'h5 == io_in_cnt ? 4'h6 : _GEN_28; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_5 = 3'h5 == io_in_cnt ? 4'h1 : _GEN_34; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_6 = 3'h5 == io_in_cnt ? 4'hc : _GEN_40; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_7 = 3'h5 == io_in_cnt ? 4'h7 : _GEN_46; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_8 = 3'h5 == io_in_cnt ? 4'h2 : _GEN_52; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_9 = 3'h5 == io_in_cnt ? 4'hd : _GEN_58; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_10 = 3'h5 == io_in_cnt ? 4'h8 : _GEN_64; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_11 = 3'h5 == io_in_cnt ? 4'h3 : _GEN_70; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_12 = 3'h5 == io_in_cnt ? 4'he : _GEN_76; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_13 = 3'h5 == io_in_cnt ? 4'h9 : _GEN_82; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_14 = 3'h5 == io_in_cnt ? 4'h4 : _GEN_88; // @[FFTDesigns.scala 3273:{17,17}]
endmodule
module PermutationsWithStreaming_6(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  input         io_in_en_5,
  input         io_in_en_6,
  input         io_in_en_7,
  input         io_in_en_8,
  input         io_in_en_9,
  input         io_in_en_10,
  input         io_in_en_11,
  input         io_in_en_12,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2634:24]
  wire [3:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2634:24]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2634:24]
  wire  RAM_Block_16_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_16_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_16_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_16_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_17_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_17_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_17_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_18_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_18_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_18_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_19_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_19_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_19_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_20_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_20_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_20_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_21_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_21_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_21_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_22_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_22_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_22_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_23_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_23_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_23_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_24_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_24_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_24_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_24_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_25_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_25_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_25_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_25_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_26_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_26_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_26_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_26_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_27_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_27_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_27_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_27_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_28_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_28_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_28_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_28_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_29_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_29_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_29_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_29_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_30_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_30_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_30_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_30_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_clock; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_31_io_in_raddr; // @[FFTDesigns.scala 2638:24]
  wire [3:0] RAM_Block_31_io_in_waddr; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_in_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_in_data_Im; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_re; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_wr; // @[FFTDesigns.scala 2638:24]
  wire  RAM_Block_31_io_en; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_out_data_Re; // @[FFTDesigns.scala 2638:24]
  wire [31:0] RAM_Block_31_io_out_data_Im; // @[FFTDesigns.scala 2638:24]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_8_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_8_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_9_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_9_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_10_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_10_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_11_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_11_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_12_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_12_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_13_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_13_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_14_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_14_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_15_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_in_15_Im; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_7; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_8; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_9; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_10; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_11; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_12; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_13; // @[FFTDesigns.scala 2641:26]
  wire [3:0] PermutationModuleStreamed_io_in_config_14; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2641:26]
  wire [31:0] PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2641:26]
  wire [2:0] M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_8; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_9; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_10; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_11; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_12; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_13; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_14; // @[FFTDesigns.scala 2642:27]
  wire [3:0] M0_Config_ROM_io_out_15; // @[FFTDesigns.scala 2642:27]
  wire [2:0] M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_8; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_9; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_10; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_11; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_12; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_13; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_14; // @[FFTDesigns.scala 2643:27]
  wire [3:0] M1_Config_ROM_io_out_15; // @[FFTDesigns.scala 2643:27]
  wire [2:0] Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2644:29]
  wire [3:0] Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2644:29]
  reg  offset_switch; // @[FFTDesigns.scala 2627:28]
  wire [5:0] lo = {io_in_en_5,io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2628:19]
  wire [12:0] _T = {io_in_en_12,io_in_en_11,io_in_en_10,io_in_en_9,io_in_en_8,io_in_en_7,io_in_en_6,lo}; // @[FFTDesigns.scala 2628:19]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2628:26]
  reg [2:0] cnt; // @[FFTDesigns.scala 2645:22]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2649:26]
  wire [2:0] _cnt_T_1 = cnt + 3'h1; // @[FFTDesigns.scala 2651:20]
  wire  _GEN_2 = cnt == 3'h5 ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2647:32 2649:23 2652:23]
  wire [3:0] _T_6 = 3'h6 * _offset_switch_T; // @[FFTDesigns.scala 2661:54]
  wire [3:0] _T_8 = M0_Config_ROM_io_out_0 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_9 = 3'h6 * offset_switch; // @[FFTDesigns.scala 2662:41]
  wire [3:0] _GEN_214 = {{1'd0}, cnt}; // @[FFTDesigns.scala 2662:31]
  wire [3:0] _T_11 = _GEN_214 + _T_9; // @[FFTDesigns.scala 2662:31]
  wire [3:0] _T_15 = _GEN_214 + _T_6; // @[FFTDesigns.scala 2664:31]
  wire [3:0] _T_18 = M1_Config_ROM_io_out_0 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_22 = M0_Config_ROM_io_out_1 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_32 = M1_Config_ROM_io_out_1 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_36 = M0_Config_ROM_io_out_2 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_46 = M1_Config_ROM_io_out_2 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_50 = M0_Config_ROM_io_out_3 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_60 = M1_Config_ROM_io_out_3 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_64 = M0_Config_ROM_io_out_4 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_74 = M1_Config_ROM_io_out_4 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_78 = M0_Config_ROM_io_out_5 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_88 = M1_Config_ROM_io_out_5 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_92 = M0_Config_ROM_io_out_6 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_102 = M1_Config_ROM_io_out_6 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_106 = M0_Config_ROM_io_out_7 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_116 = M1_Config_ROM_io_out_7 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_120 = M0_Config_ROM_io_out_8 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_130 = M1_Config_ROM_io_out_8 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_134 = M0_Config_ROM_io_out_9 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_144 = M1_Config_ROM_io_out_9 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_148 = M0_Config_ROM_io_out_10 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_158 = M1_Config_ROM_io_out_10 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_162 = M0_Config_ROM_io_out_11 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_172 = M1_Config_ROM_io_out_11 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_176 = M0_Config_ROM_io_out_12 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_186 = M1_Config_ROM_io_out_12 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_190 = M0_Config_ROM_io_out_13 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_200 = M1_Config_ROM_io_out_13 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_204 = M0_Config_ROM_io_out_14 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_214 = M1_Config_ROM_io_out_14 + _T_9; // @[FFTDesigns.scala 2665:44]
  wire [3:0] _T_218 = M0_Config_ROM_io_out_15 + _T_6; // @[FFTDesigns.scala 2661:44]
  wire [3:0] _T_228 = M1_Config_ROM_io_out_15 + _T_9; // @[FFTDesigns.scala 2665:44]
  RAM_Block_192 RAM_Block ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_1 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_2 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_3 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_4 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_5 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_6 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_7 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_8 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_9 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_10 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_11 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_12 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_13 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_14 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_15 ( // @[FFTDesigns.scala 2634:24]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_16 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_16_clock),
    .io_in_raddr(RAM_Block_16_io_in_raddr),
    .io_in_waddr(RAM_Block_16_io_in_waddr),
    .io_in_data_Re(RAM_Block_16_io_in_data_Re),
    .io_in_data_Im(RAM_Block_16_io_in_data_Im),
    .io_re(RAM_Block_16_io_re),
    .io_wr(RAM_Block_16_io_wr),
    .io_en(RAM_Block_16_io_en),
    .io_out_data_Re(RAM_Block_16_io_out_data_Re),
    .io_out_data_Im(RAM_Block_16_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_17 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_17_clock),
    .io_in_raddr(RAM_Block_17_io_in_raddr),
    .io_in_waddr(RAM_Block_17_io_in_waddr),
    .io_in_data_Re(RAM_Block_17_io_in_data_Re),
    .io_in_data_Im(RAM_Block_17_io_in_data_Im),
    .io_re(RAM_Block_17_io_re),
    .io_wr(RAM_Block_17_io_wr),
    .io_en(RAM_Block_17_io_en),
    .io_out_data_Re(RAM_Block_17_io_out_data_Re),
    .io_out_data_Im(RAM_Block_17_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_18 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_18_clock),
    .io_in_raddr(RAM_Block_18_io_in_raddr),
    .io_in_waddr(RAM_Block_18_io_in_waddr),
    .io_in_data_Re(RAM_Block_18_io_in_data_Re),
    .io_in_data_Im(RAM_Block_18_io_in_data_Im),
    .io_re(RAM_Block_18_io_re),
    .io_wr(RAM_Block_18_io_wr),
    .io_en(RAM_Block_18_io_en),
    .io_out_data_Re(RAM_Block_18_io_out_data_Re),
    .io_out_data_Im(RAM_Block_18_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_19 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_19_clock),
    .io_in_raddr(RAM_Block_19_io_in_raddr),
    .io_in_waddr(RAM_Block_19_io_in_waddr),
    .io_in_data_Re(RAM_Block_19_io_in_data_Re),
    .io_in_data_Im(RAM_Block_19_io_in_data_Im),
    .io_re(RAM_Block_19_io_re),
    .io_wr(RAM_Block_19_io_wr),
    .io_en(RAM_Block_19_io_en),
    .io_out_data_Re(RAM_Block_19_io_out_data_Re),
    .io_out_data_Im(RAM_Block_19_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_20 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_20_clock),
    .io_in_raddr(RAM_Block_20_io_in_raddr),
    .io_in_waddr(RAM_Block_20_io_in_waddr),
    .io_in_data_Re(RAM_Block_20_io_in_data_Re),
    .io_in_data_Im(RAM_Block_20_io_in_data_Im),
    .io_re(RAM_Block_20_io_re),
    .io_wr(RAM_Block_20_io_wr),
    .io_en(RAM_Block_20_io_en),
    .io_out_data_Re(RAM_Block_20_io_out_data_Re),
    .io_out_data_Im(RAM_Block_20_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_21 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_21_clock),
    .io_in_raddr(RAM_Block_21_io_in_raddr),
    .io_in_waddr(RAM_Block_21_io_in_waddr),
    .io_in_data_Re(RAM_Block_21_io_in_data_Re),
    .io_in_data_Im(RAM_Block_21_io_in_data_Im),
    .io_re(RAM_Block_21_io_re),
    .io_wr(RAM_Block_21_io_wr),
    .io_en(RAM_Block_21_io_en),
    .io_out_data_Re(RAM_Block_21_io_out_data_Re),
    .io_out_data_Im(RAM_Block_21_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_22 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_22_clock),
    .io_in_raddr(RAM_Block_22_io_in_raddr),
    .io_in_waddr(RAM_Block_22_io_in_waddr),
    .io_in_data_Re(RAM_Block_22_io_in_data_Re),
    .io_in_data_Im(RAM_Block_22_io_in_data_Im),
    .io_re(RAM_Block_22_io_re),
    .io_wr(RAM_Block_22_io_wr),
    .io_en(RAM_Block_22_io_en),
    .io_out_data_Re(RAM_Block_22_io_out_data_Re),
    .io_out_data_Im(RAM_Block_22_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_23 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_23_clock),
    .io_in_raddr(RAM_Block_23_io_in_raddr),
    .io_in_waddr(RAM_Block_23_io_in_waddr),
    .io_in_data_Re(RAM_Block_23_io_in_data_Re),
    .io_in_data_Im(RAM_Block_23_io_in_data_Im),
    .io_re(RAM_Block_23_io_re),
    .io_wr(RAM_Block_23_io_wr),
    .io_en(RAM_Block_23_io_en),
    .io_out_data_Re(RAM_Block_23_io_out_data_Re),
    .io_out_data_Im(RAM_Block_23_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_24 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_24_clock),
    .io_in_raddr(RAM_Block_24_io_in_raddr),
    .io_in_waddr(RAM_Block_24_io_in_waddr),
    .io_in_data_Re(RAM_Block_24_io_in_data_Re),
    .io_in_data_Im(RAM_Block_24_io_in_data_Im),
    .io_re(RAM_Block_24_io_re),
    .io_wr(RAM_Block_24_io_wr),
    .io_en(RAM_Block_24_io_en),
    .io_out_data_Re(RAM_Block_24_io_out_data_Re),
    .io_out_data_Im(RAM_Block_24_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_25 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_25_clock),
    .io_in_raddr(RAM_Block_25_io_in_raddr),
    .io_in_waddr(RAM_Block_25_io_in_waddr),
    .io_in_data_Re(RAM_Block_25_io_in_data_Re),
    .io_in_data_Im(RAM_Block_25_io_in_data_Im),
    .io_re(RAM_Block_25_io_re),
    .io_wr(RAM_Block_25_io_wr),
    .io_en(RAM_Block_25_io_en),
    .io_out_data_Re(RAM_Block_25_io_out_data_Re),
    .io_out_data_Im(RAM_Block_25_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_26 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_26_clock),
    .io_in_raddr(RAM_Block_26_io_in_raddr),
    .io_in_waddr(RAM_Block_26_io_in_waddr),
    .io_in_data_Re(RAM_Block_26_io_in_data_Re),
    .io_in_data_Im(RAM_Block_26_io_in_data_Im),
    .io_re(RAM_Block_26_io_re),
    .io_wr(RAM_Block_26_io_wr),
    .io_en(RAM_Block_26_io_en),
    .io_out_data_Re(RAM_Block_26_io_out_data_Re),
    .io_out_data_Im(RAM_Block_26_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_27 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_27_clock),
    .io_in_raddr(RAM_Block_27_io_in_raddr),
    .io_in_waddr(RAM_Block_27_io_in_waddr),
    .io_in_data_Re(RAM_Block_27_io_in_data_Re),
    .io_in_data_Im(RAM_Block_27_io_in_data_Im),
    .io_re(RAM_Block_27_io_re),
    .io_wr(RAM_Block_27_io_wr),
    .io_en(RAM_Block_27_io_en),
    .io_out_data_Re(RAM_Block_27_io_out_data_Re),
    .io_out_data_Im(RAM_Block_27_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_28 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_28_clock),
    .io_in_raddr(RAM_Block_28_io_in_raddr),
    .io_in_waddr(RAM_Block_28_io_in_waddr),
    .io_in_data_Re(RAM_Block_28_io_in_data_Re),
    .io_in_data_Im(RAM_Block_28_io_in_data_Im),
    .io_re(RAM_Block_28_io_re),
    .io_wr(RAM_Block_28_io_wr),
    .io_en(RAM_Block_28_io_en),
    .io_out_data_Re(RAM_Block_28_io_out_data_Re),
    .io_out_data_Im(RAM_Block_28_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_29 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_29_clock),
    .io_in_raddr(RAM_Block_29_io_in_raddr),
    .io_in_waddr(RAM_Block_29_io_in_waddr),
    .io_in_data_Re(RAM_Block_29_io_in_data_Re),
    .io_in_data_Im(RAM_Block_29_io_in_data_Im),
    .io_re(RAM_Block_29_io_re),
    .io_wr(RAM_Block_29_io_wr),
    .io_en(RAM_Block_29_io_en),
    .io_out_data_Re(RAM_Block_29_io_out_data_Re),
    .io_out_data_Im(RAM_Block_29_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_30 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_30_clock),
    .io_in_raddr(RAM_Block_30_io_in_raddr),
    .io_in_waddr(RAM_Block_30_io_in_waddr),
    .io_in_data_Re(RAM_Block_30_io_in_data_Re),
    .io_in_data_Im(RAM_Block_30_io_in_data_Im),
    .io_re(RAM_Block_30_io_re),
    .io_wr(RAM_Block_30_io_wr),
    .io_en(RAM_Block_30_io_en),
    .io_out_data_Re(RAM_Block_30_io_out_data_Re),
    .io_out_data_Im(RAM_Block_30_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_31 ( // @[FFTDesigns.scala 2638:24]
    .clock(RAM_Block_31_clock),
    .io_in_raddr(RAM_Block_31_io_in_raddr),
    .io_in_waddr(RAM_Block_31_io_in_waddr),
    .io_in_data_Re(RAM_Block_31_io_in_data_Re),
    .io_in_data_Im(RAM_Block_31_io_in_data_Im),
    .io_re(RAM_Block_31_io_re),
    .io_wr(RAM_Block_31_io_wr),
    .io_en(RAM_Block_31_io_en),
    .io_out_data_Re(RAM_Block_31_io_out_data_Re),
    .io_out_data_Im(RAM_Block_31_io_out_data_Im)
  );
  PermutationModuleStreamed PermutationModuleStreamed ( // @[FFTDesigns.scala 2641:26]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_8_Re(PermutationModuleStreamed_io_in_8_Re),
    .io_in_8_Im(PermutationModuleStreamed_io_in_8_Im),
    .io_in_9_Re(PermutationModuleStreamed_io_in_9_Re),
    .io_in_9_Im(PermutationModuleStreamed_io_in_9_Im),
    .io_in_10_Re(PermutationModuleStreamed_io_in_10_Re),
    .io_in_10_Im(PermutationModuleStreamed_io_in_10_Im),
    .io_in_11_Re(PermutationModuleStreamed_io_in_11_Re),
    .io_in_11_Im(PermutationModuleStreamed_io_in_11_Im),
    .io_in_12_Re(PermutationModuleStreamed_io_in_12_Re),
    .io_in_12_Im(PermutationModuleStreamed_io_in_12_Im),
    .io_in_13_Re(PermutationModuleStreamed_io_in_13_Re),
    .io_in_13_Im(PermutationModuleStreamed_io_in_13_Im),
    .io_in_14_Re(PermutationModuleStreamed_io_in_14_Re),
    .io_in_14_Im(PermutationModuleStreamed_io_in_14_Im),
    .io_in_15_Re(PermutationModuleStreamed_io_in_15_Re),
    .io_in_15_Im(PermutationModuleStreamed_io_in_15_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_in_config_7(PermutationModuleStreamed_io_in_config_7),
    .io_in_config_8(PermutationModuleStreamed_io_in_config_8),
    .io_in_config_9(PermutationModuleStreamed_io_in_config_9),
    .io_in_config_10(PermutationModuleStreamed_io_in_config_10),
    .io_in_config_11(PermutationModuleStreamed_io_in_config_11),
    .io_in_config_12(PermutationModuleStreamed_io_in_config_12),
    .io_in_config_13(PermutationModuleStreamed_io_in_config_13),
    .io_in_config_14(PermutationModuleStreamed_io_in_config_14),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im),
    .io_out_8_Re(PermutationModuleStreamed_io_out_8_Re),
    .io_out_8_Im(PermutationModuleStreamed_io_out_8_Im),
    .io_out_9_Re(PermutationModuleStreamed_io_out_9_Re),
    .io_out_9_Im(PermutationModuleStreamed_io_out_9_Im),
    .io_out_10_Re(PermutationModuleStreamed_io_out_10_Re),
    .io_out_10_Im(PermutationModuleStreamed_io_out_10_Im),
    .io_out_11_Re(PermutationModuleStreamed_io_out_11_Re),
    .io_out_11_Im(PermutationModuleStreamed_io_out_11_Im),
    .io_out_12_Re(PermutationModuleStreamed_io_out_12_Re),
    .io_out_12_Im(PermutationModuleStreamed_io_out_12_Im),
    .io_out_13_Re(PermutationModuleStreamed_io_out_13_Re),
    .io_out_13_Im(PermutationModuleStreamed_io_out_13_Im),
    .io_out_14_Re(PermutationModuleStreamed_io_out_14_Re),
    .io_out_14_Im(PermutationModuleStreamed_io_out_14_Im),
    .io_out_15_Re(PermutationModuleStreamed_io_out_15_Re),
    .io_out_15_Im(PermutationModuleStreamed_io_out_15_Im)
  );
  M0_Config_ROM_6 M0_Config_ROM ( // @[FFTDesigns.scala 2642:27]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7),
    .io_out_8(M0_Config_ROM_io_out_8),
    .io_out_9(M0_Config_ROM_io_out_9),
    .io_out_10(M0_Config_ROM_io_out_10),
    .io_out_11(M0_Config_ROM_io_out_11),
    .io_out_12(M0_Config_ROM_io_out_12),
    .io_out_13(M0_Config_ROM_io_out_13),
    .io_out_14(M0_Config_ROM_io_out_14),
    .io_out_15(M0_Config_ROM_io_out_15)
  );
  M1_Config_ROM_6 M1_Config_ROM ( // @[FFTDesigns.scala 2643:27]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7),
    .io_out_8(M1_Config_ROM_io_out_8),
    .io_out_9(M1_Config_ROM_io_out_9),
    .io_out_10(M1_Config_ROM_io_out_10),
    .io_out_11(M1_Config_ROM_io_out_11),
    .io_out_12(M1_Config_ROM_io_out_12),
    .io_out_13(M1_Config_ROM_io_out_13),
    .io_out_14(M1_Config_ROM_io_out_14),
    .io_out_15(M1_Config_ROM_io_out_15)
  );
  Streaming_Permute_Config_6 Streaming_Permute_Config ( // @[FFTDesigns.scala 2644:29]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6),
    .io_out_7(Streaming_Permute_Config_io_out_7),
    .io_out_8(Streaming_Permute_Config_io_out_8),
    .io_out_9(Streaming_Permute_Config_io_out_9),
    .io_out_10(Streaming_Permute_Config_io_out_10),
    .io_out_11(Streaming_Permute_Config_io_out_11),
    .io_out_12(Streaming_Permute_Config_io_out_12),
    .io_out_13(Streaming_Permute_Config_io_out_13),
    .io_out_14(Streaming_Permute_Config_io_out_14)
  );
  assign io_out_0_Re = RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_0_Im = RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Re = RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_1_Im = RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Re = RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_2_Im = RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Re = RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_3_Im = RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Re = RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_4_Im = RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Re = RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_5_Im = RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Re = RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_6_Im = RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Re = RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_7_Im = RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_8_Re = RAM_Block_24_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_8_Im = RAM_Block_24_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_9_Re = RAM_Block_25_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_9_Im = RAM_Block_25_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_10_Re = RAM_Block_26_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_10_Im = RAM_Block_26_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_11_Re = RAM_Block_27_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_11_Im = RAM_Block_27_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_12_Re = RAM_Block_28_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_12_Im = RAM_Block_28_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_13_Re = RAM_Block_29_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_13_Im = RAM_Block_29_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_14_Re = RAM_Block_30_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_14_Im = RAM_Block_30_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_15_Re = RAM_Block_31_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign io_out_15_Im = RAM_Block_31_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2670:19 2689:19]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = _T_1 ? _T_8 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_io_in_data_Re = io_in_0_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_in_data_Im = io_in_0_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = _T_1 ? _T_22 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_1_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_1_io_in_data_Re = io_in_1_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_in_data_Im = io_in_1_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = _T_1 ? _T_36 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_2_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_2_io_in_data_Re = io_in_2_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_in_data_Im = io_in_2_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = _T_1 ? _T_50 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_3_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_3_io_in_data_Re = io_in_3_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_in_data_Im = io_in_3_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = _T_1 ? _T_64 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_4_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_4_io_in_data_Re = io_in_4_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_in_data_Im = io_in_4_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = _T_1 ? _T_78 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_5_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_5_io_in_data_Re = io_in_5_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_in_data_Im = io_in_5_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = _T_1 ? _T_92 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_6_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_6_io_in_data_Re = io_in_6_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_in_data_Im = io_in_6_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = _T_1 ? _T_106 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_7_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_7_io_in_data_Re = io_in_7_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_in_data_Im = io_in_7_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = _T_1 ? _T_120 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_8_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_8_io_in_data_Re = io_in_8_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_8_io_in_data_Im = io_in_8_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = _T_1 ? _T_134 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_9_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_9_io_in_data_Re = io_in_9_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_9_io_in_data_Im = io_in_9_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = _T_1 ? _T_148 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_10_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_10_io_in_data_Re = io_in_10_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_10_io_in_data_Im = io_in_10_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = _T_1 ? _T_162 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_11_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_11_io_in_data_Re = io_in_11_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_11_io_in_data_Im = io_in_11_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = _T_1 ? _T_176 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_12_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_12_io_in_data_Re = io_in_12_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_12_io_in_data_Im = io_in_12_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = _T_1 ? _T_190 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_13_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_13_io_in_data_Re = io_in_13_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_13_io_in_data_Im = io_in_13_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = _T_1 ? _T_204 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_14_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_14_io_in_data_Re = io_in_14_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_14_io_in_data_Im = io_in_14_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = _T_1 ? _T_218 : 4'h0; // @[FFTDesigns.scala 2646:30 2661:24 2680:24]
  assign RAM_Block_15_io_in_waddr = _T_1 ? _T_11 : 4'h0; // @[FFTDesigns.scala 2646:30 2662:24 2681:24]
  assign RAM_Block_15_io_in_data_Re = io_in_15_Re; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_15_io_in_data_Im = io_in_15_Im; // @[FFTDesigns.scala 2646:30 2663:23 2682:23]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_clock = clock;
  assign RAM_Block_16_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_16_io_in_waddr = _T_1 ? _T_18 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_16_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_16_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_16_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_16_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_clock = clock;
  assign RAM_Block_17_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_17_io_in_waddr = _T_1 ? _T_32 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_17_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_17_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_17_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_17_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_clock = clock;
  assign RAM_Block_18_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_18_io_in_waddr = _T_1 ? _T_46 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_18_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_18_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_18_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_18_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_clock = clock;
  assign RAM_Block_19_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_19_io_in_waddr = _T_1 ? _T_60 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_19_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_19_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_19_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_19_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_clock = clock;
  assign RAM_Block_20_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_20_io_in_waddr = _T_1 ? _T_74 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_20_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_20_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_20_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_20_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_clock = clock;
  assign RAM_Block_21_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_21_io_in_waddr = _T_1 ? _T_88 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_21_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_21_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_21_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_21_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_clock = clock;
  assign RAM_Block_22_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_22_io_in_waddr = _T_1 ? _T_102 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_22_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_22_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_22_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_22_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_clock = clock;
  assign RAM_Block_23_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_23_io_in_waddr = _T_1 ? _T_116 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_23_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_23_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_23_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_23_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_clock = clock;
  assign RAM_Block_24_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_24_io_in_waddr = _T_1 ? _T_130 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_24_io_in_data_Re = PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_24_io_in_data_Im = PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_24_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_24_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_clock = clock;
  assign RAM_Block_25_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_25_io_in_waddr = _T_1 ? _T_144 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_25_io_in_data_Re = PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_25_io_in_data_Im = PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_25_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_25_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_clock = clock;
  assign RAM_Block_26_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_26_io_in_waddr = _T_1 ? _T_158 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_26_io_in_data_Re = PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_26_io_in_data_Im = PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_26_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_26_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_clock = clock;
  assign RAM_Block_27_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_27_io_in_waddr = _T_1 ? _T_172 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_27_io_in_data_Re = PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_27_io_in_data_Im = PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_27_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_27_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_clock = clock;
  assign RAM_Block_28_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_28_io_in_waddr = _T_1 ? _T_186 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_28_io_in_data_Re = PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_28_io_in_data_Im = PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_28_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_28_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_clock = clock;
  assign RAM_Block_29_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_29_io_in_waddr = _T_1 ? _T_200 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_29_io_in_data_Re = PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_29_io_in_data_Im = PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_29_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_29_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_clock = clock;
  assign RAM_Block_30_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_30_io_in_waddr = _T_1 ? _T_214 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_30_io_in_data_Re = PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_30_io_in_data_Im = PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_30_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_30_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_clock = clock;
  assign RAM_Block_31_io_in_raddr = _T_1 ? _T_15 : 4'h0; // @[FFTDesigns.scala 2646:30 2664:24 2683:24]
  assign RAM_Block_31_io_in_waddr = _T_1 ? _T_228 : 4'h0; // @[FFTDesigns.scala 2646:30 2665:24 2684:24]
  assign RAM_Block_31_io_in_data_Re = PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_31_io_in_data_Im = PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2646:30 2666:23 2685:23]
  assign RAM_Block_31_io_re = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_io_wr = |_T; // @[FFTDesigns.scala 2646:26]
  assign RAM_Block_31_io_en = |_T; // @[FFTDesigns.scala 2646:26]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_8_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_8_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_9_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_9_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_10_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_10_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_11_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_11_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_12_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_12_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_13_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_13_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_14_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_14_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_15_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_15_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2646:30 2668:24 2687:24]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_7 = Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_8 = Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_9 = Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_10 = Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_11 = Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_12 = Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_13 = Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign PermutationModuleStreamed_io_in_config_14 = Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2646:30 2667:31 2686:31]
  assign M0_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2694:22]
  assign M1_Config_ROM_io_in_cnt = cnt; // @[FFTDesigns.scala 2695:22]
  assign Streaming_Permute_Config_io_in_cnt = cnt; // @[FFTDesigns.scala 2696:24]
  always @(posedge clock) begin
    offset_switch <= _T_1 & _GEN_2; // @[FFTDesigns.scala 2646:30 2691:21]
    if (reset) begin // @[FFTDesigns.scala 2645:22]
      cnt <= 3'h0; // @[FFTDesigns.scala 2645:22]
    end else if (_T_1) begin // @[FFTDesigns.scala 2646:30]
      if (cnt == 3'h5) begin // @[FFTDesigns.scala 2647:32]
        cnt <= 3'h0; // @[FFTDesigns.scala 2648:13]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2651:13]
      end
    end else begin
      cnt <= 3'h0; // @[FFTDesigns.scala 2692:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_Block_224(
  input         clock,
  input  [2:0]  io_in_raddr,
  input  [2:0]  io_in_waddr,
  input  [31:0] io_in_data_Re,
  input  [31:0] io_in_data_Im,
  input         io_re,
  input         io_wr,
  input         io_en,
  output [31:0] io_out_data_Re,
  output [31:0] io_out_data_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_0_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_1_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_2_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_3_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_4_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_5_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_6_Im; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Re; // @[FFTDesigns.scala 3286:18]
  reg [31:0] mem_7_Im; // @[FFTDesigns.scala 3286:18]
  wire [31:0] _GEN_33 = 3'h1 == io_in_raddr ? mem_1_Im : mem_0_Im; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_34 = 3'h2 == io_in_raddr ? mem_2_Im : _GEN_33; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_35 = 3'h3 == io_in_raddr ? mem_3_Im : _GEN_34; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_36 = 3'h4 == io_in_raddr ? mem_4_Im : _GEN_35; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_37 = 3'h5 == io_in_raddr ? mem_5_Im : _GEN_36; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_38 = 3'h6 == io_in_raddr ? mem_6_Im : _GEN_37; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_39 = 3'h7 == io_in_raddr ? mem_7_Im : _GEN_38; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_41 = 3'h1 == io_in_raddr ? mem_1_Re : mem_0_Re; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_42 = 3'h2 == io_in_raddr ? mem_2_Re : _GEN_41; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_43 = 3'h3 == io_in_raddr ? mem_3_Re : _GEN_42; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_44 = 3'h4 == io_in_raddr ? mem_4_Re : _GEN_43; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_45 = 3'h5 == io_in_raddr ? mem_5_Re : _GEN_44; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_46 = 3'h6 == io_in_raddr ? mem_6_Re : _GEN_45; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_47 = 3'h7 == io_in_raddr ? mem_7_Re : _GEN_46; // @[FFTDesigns.scala 3292:{21,21}]
  wire [31:0] _GEN_48 = io_re ? _GEN_39 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3295:24]
  wire [31:0] _GEN_49 = io_re ? _GEN_47 : 32'h0; // @[FFTDesigns.scala 3291:18 3292:21 3294:24]
  assign io_out_data_Re = io_en ? _GEN_49 : 32'h0; // @[FFTDesigns.scala 3287:16 3298:22]
  assign io_out_data_Im = io_en ? _GEN_48 : 32'h0; // @[FFTDesigns.scala 3287:16 3299:22]
  always @(posedge clock) begin
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h0 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_0_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h1 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_1_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h2 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_2_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h3 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_3_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h4 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_4_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h5 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_5_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h6 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_6_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Re <= io_in_data_Re; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3287:16]
      if (io_wr) begin // @[FFTDesigns.scala 3288:18]
        if (3'h7 == io_in_waddr) begin // @[FFTDesigns.scala 3289:26]
          mem_7_Im <= io_in_data_Im; // @[FFTDesigns.scala 3289:26]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_3_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_4_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_4_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_5_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_5_Im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_6_Re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_6_Im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_7_Re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_7_Im = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PermutationModuleStreamed_7(
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input  [4:0]  io_in_config_0,
  input  [4:0]  io_in_config_1,
  input  [4:0]  io_in_config_2,
  input  [4:0]  io_in_config_3,
  input  [4:0]  io_in_config_4,
  input  [4:0]  io_in_config_5,
  input  [4:0]  io_in_config_6,
  input  [4:0]  io_in_config_7,
  input  [4:0]  io_in_config_8,
  input  [4:0]  io_in_config_9,
  input  [4:0]  io_in_config_10,
  input  [4:0]  io_in_config_11,
  input  [4:0]  io_in_config_12,
  input  [4:0]  io_in_config_13,
  input  [4:0]  io_in_config_14,
  input  [4:0]  io_in_config_15,
  input  [4:0]  io_in_config_16,
  input  [4:0]  io_in_config_17,
  input  [4:0]  io_in_config_18,
  input  [4:0]  io_in_config_19,
  input  [4:0]  io_in_config_20,
  input  [4:0]  io_in_config_21,
  input  [4:0]  io_in_config_22,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im
);
  wire  _T = io_in_config_0 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_1 = io_in_config_1 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_2 = io_in_config_2 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_3 = io_in_config_3 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_4 = io_in_config_4 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_5 = io_in_config_5 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_6 = io_in_config_6 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_7 = io_in_config_7 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_8 = io_in_config_8 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_9 = io_in_config_9 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_10 = io_in_config_10 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_11 = io_in_config_11 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_12 = io_in_config_12 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_13 = io_in_config_13 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_14 = io_in_config_14 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_15 = io_in_config_15 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_16 = io_in_config_16 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_17 = io_in_config_17 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_18 = io_in_config_18 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_19 = io_in_config_19 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_20 = io_in_config_20 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_21 = io_in_config_21 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_22 = io_in_config_22 == 5'h0; // @[FFTDesigns.scala 3194:35]
  wire  _T_24 = io_in_config_0 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_25 = io_in_config_1 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_26 = io_in_config_2 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_27 = io_in_config_3 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_28 = io_in_config_4 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_29 = io_in_config_5 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_30 = io_in_config_6 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_31 = io_in_config_7 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_32 = io_in_config_8 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_33 = io_in_config_9 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_34 = io_in_config_10 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_35 = io_in_config_11 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_36 = io_in_config_12 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_37 = io_in_config_13 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_38 = io_in_config_14 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_39 = io_in_config_15 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_40 = io_in_config_16 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_41 = io_in_config_17 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_42 = io_in_config_18 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_43 = io_in_config_19 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_44 = io_in_config_20 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_45 = io_in_config_21 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_46 = io_in_config_22 == 5'h1; // @[FFTDesigns.scala 3194:35]
  wire  _T_48 = io_in_config_0 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_49 = io_in_config_1 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_50 = io_in_config_2 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_51 = io_in_config_3 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_52 = io_in_config_4 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_53 = io_in_config_5 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_54 = io_in_config_6 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_55 = io_in_config_7 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_56 = io_in_config_8 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_57 = io_in_config_9 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_58 = io_in_config_10 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_59 = io_in_config_11 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_60 = io_in_config_12 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_61 = io_in_config_13 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_62 = io_in_config_14 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_63 = io_in_config_15 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_64 = io_in_config_16 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_65 = io_in_config_17 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_66 = io_in_config_18 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_67 = io_in_config_19 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_68 = io_in_config_20 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_69 = io_in_config_21 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_70 = io_in_config_22 == 5'h2; // @[FFTDesigns.scala 3194:35]
  wire  _T_72 = io_in_config_0 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_73 = io_in_config_1 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_74 = io_in_config_2 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_75 = io_in_config_3 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_76 = io_in_config_4 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_77 = io_in_config_5 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_78 = io_in_config_6 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_79 = io_in_config_7 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_80 = io_in_config_8 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_81 = io_in_config_9 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_82 = io_in_config_10 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_83 = io_in_config_11 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_84 = io_in_config_12 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_85 = io_in_config_13 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_86 = io_in_config_14 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_87 = io_in_config_15 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_88 = io_in_config_16 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_89 = io_in_config_17 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_90 = io_in_config_18 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_91 = io_in_config_19 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_92 = io_in_config_20 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_93 = io_in_config_21 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_94 = io_in_config_22 == 5'h3; // @[FFTDesigns.scala 3194:35]
  wire  _T_96 = io_in_config_0 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_97 = io_in_config_1 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_98 = io_in_config_2 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_99 = io_in_config_3 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_100 = io_in_config_4 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_101 = io_in_config_5 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_102 = io_in_config_6 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_103 = io_in_config_7 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_104 = io_in_config_8 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_105 = io_in_config_9 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_106 = io_in_config_10 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_107 = io_in_config_11 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_108 = io_in_config_12 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_109 = io_in_config_13 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_110 = io_in_config_14 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_111 = io_in_config_15 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_112 = io_in_config_16 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_113 = io_in_config_17 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_114 = io_in_config_18 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_115 = io_in_config_19 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_116 = io_in_config_20 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_117 = io_in_config_21 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_118 = io_in_config_22 == 5'h4; // @[FFTDesigns.scala 3194:35]
  wire  _T_120 = io_in_config_0 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_121 = io_in_config_1 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_122 = io_in_config_2 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_123 = io_in_config_3 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_124 = io_in_config_4 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_125 = io_in_config_5 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_126 = io_in_config_6 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_127 = io_in_config_7 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_128 = io_in_config_8 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_129 = io_in_config_9 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_130 = io_in_config_10 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_131 = io_in_config_11 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_132 = io_in_config_12 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_133 = io_in_config_13 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_134 = io_in_config_14 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_135 = io_in_config_15 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_136 = io_in_config_16 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_137 = io_in_config_17 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_138 = io_in_config_18 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_139 = io_in_config_19 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_140 = io_in_config_20 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_141 = io_in_config_21 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_142 = io_in_config_22 == 5'h5; // @[FFTDesigns.scala 3194:35]
  wire  _T_144 = io_in_config_0 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_145 = io_in_config_1 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_146 = io_in_config_2 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_147 = io_in_config_3 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_148 = io_in_config_4 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_149 = io_in_config_5 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_150 = io_in_config_6 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_151 = io_in_config_7 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_152 = io_in_config_8 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_153 = io_in_config_9 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_154 = io_in_config_10 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_155 = io_in_config_11 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_156 = io_in_config_12 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_157 = io_in_config_13 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_158 = io_in_config_14 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_159 = io_in_config_15 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_160 = io_in_config_16 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_161 = io_in_config_17 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_162 = io_in_config_18 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_163 = io_in_config_19 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_164 = io_in_config_20 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_165 = io_in_config_21 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_166 = io_in_config_22 == 5'h6; // @[FFTDesigns.scala 3194:35]
  wire  _T_168 = io_in_config_0 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_169 = io_in_config_1 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_170 = io_in_config_2 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_171 = io_in_config_3 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_172 = io_in_config_4 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_173 = io_in_config_5 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_174 = io_in_config_6 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_175 = io_in_config_7 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_176 = io_in_config_8 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_177 = io_in_config_9 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_178 = io_in_config_10 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_179 = io_in_config_11 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_180 = io_in_config_12 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_181 = io_in_config_13 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_182 = io_in_config_14 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_183 = io_in_config_15 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_184 = io_in_config_16 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_185 = io_in_config_17 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_186 = io_in_config_18 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_187 = io_in_config_19 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_188 = io_in_config_20 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_189 = io_in_config_21 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_190 = io_in_config_22 == 5'h7; // @[FFTDesigns.scala 3194:35]
  wire  _T_192 = io_in_config_0 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_193 = io_in_config_1 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_194 = io_in_config_2 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_195 = io_in_config_3 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_196 = io_in_config_4 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_197 = io_in_config_5 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_198 = io_in_config_6 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_199 = io_in_config_7 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_200 = io_in_config_8 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_201 = io_in_config_9 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_202 = io_in_config_10 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_203 = io_in_config_11 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_204 = io_in_config_12 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_205 = io_in_config_13 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_206 = io_in_config_14 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_207 = io_in_config_15 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_208 = io_in_config_16 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_209 = io_in_config_17 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_210 = io_in_config_18 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_211 = io_in_config_19 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_212 = io_in_config_20 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_213 = io_in_config_21 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_214 = io_in_config_22 == 5'h8; // @[FFTDesigns.scala 3194:35]
  wire  _T_216 = io_in_config_0 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_217 = io_in_config_1 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_218 = io_in_config_2 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_219 = io_in_config_3 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_220 = io_in_config_4 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_221 = io_in_config_5 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_222 = io_in_config_6 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_223 = io_in_config_7 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_224 = io_in_config_8 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_225 = io_in_config_9 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_226 = io_in_config_10 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_227 = io_in_config_11 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_228 = io_in_config_12 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_229 = io_in_config_13 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_230 = io_in_config_14 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_231 = io_in_config_15 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_232 = io_in_config_16 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_233 = io_in_config_17 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_234 = io_in_config_18 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_235 = io_in_config_19 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_236 = io_in_config_20 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_237 = io_in_config_21 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_238 = io_in_config_22 == 5'h9; // @[FFTDesigns.scala 3194:35]
  wire  _T_240 = io_in_config_0 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_241 = io_in_config_1 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_242 = io_in_config_2 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_243 = io_in_config_3 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_244 = io_in_config_4 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_245 = io_in_config_5 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_246 = io_in_config_6 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_247 = io_in_config_7 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_248 = io_in_config_8 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_249 = io_in_config_9 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_250 = io_in_config_10 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_251 = io_in_config_11 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_252 = io_in_config_12 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_253 = io_in_config_13 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_254 = io_in_config_14 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_255 = io_in_config_15 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_256 = io_in_config_16 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_257 = io_in_config_17 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_258 = io_in_config_18 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_259 = io_in_config_19 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_260 = io_in_config_20 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_261 = io_in_config_21 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_262 = io_in_config_22 == 5'ha; // @[FFTDesigns.scala 3194:35]
  wire  _T_264 = io_in_config_0 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_265 = io_in_config_1 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_266 = io_in_config_2 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_267 = io_in_config_3 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_268 = io_in_config_4 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_269 = io_in_config_5 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_270 = io_in_config_6 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_271 = io_in_config_7 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_272 = io_in_config_8 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_273 = io_in_config_9 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_274 = io_in_config_10 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_275 = io_in_config_11 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_276 = io_in_config_12 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_277 = io_in_config_13 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_278 = io_in_config_14 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_279 = io_in_config_15 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_280 = io_in_config_16 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_281 = io_in_config_17 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_282 = io_in_config_18 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_283 = io_in_config_19 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_284 = io_in_config_20 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_285 = io_in_config_21 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_286 = io_in_config_22 == 5'hb; // @[FFTDesigns.scala 3194:35]
  wire  _T_288 = io_in_config_0 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_289 = io_in_config_1 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_290 = io_in_config_2 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_291 = io_in_config_3 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_292 = io_in_config_4 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_293 = io_in_config_5 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_294 = io_in_config_6 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_295 = io_in_config_7 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_296 = io_in_config_8 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_297 = io_in_config_9 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_298 = io_in_config_10 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_299 = io_in_config_11 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_300 = io_in_config_12 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_301 = io_in_config_13 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_302 = io_in_config_14 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_303 = io_in_config_15 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_304 = io_in_config_16 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_305 = io_in_config_17 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_306 = io_in_config_18 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_307 = io_in_config_19 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_308 = io_in_config_20 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_309 = io_in_config_21 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_310 = io_in_config_22 == 5'hc; // @[FFTDesigns.scala 3194:35]
  wire  _T_312 = io_in_config_0 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_313 = io_in_config_1 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_314 = io_in_config_2 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_315 = io_in_config_3 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_316 = io_in_config_4 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_317 = io_in_config_5 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_318 = io_in_config_6 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_319 = io_in_config_7 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_320 = io_in_config_8 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_321 = io_in_config_9 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_322 = io_in_config_10 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_323 = io_in_config_11 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_324 = io_in_config_12 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_325 = io_in_config_13 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_326 = io_in_config_14 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_327 = io_in_config_15 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_328 = io_in_config_16 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_329 = io_in_config_17 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_330 = io_in_config_18 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_331 = io_in_config_19 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_332 = io_in_config_20 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_333 = io_in_config_21 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_334 = io_in_config_22 == 5'hd; // @[FFTDesigns.scala 3194:35]
  wire  _T_336 = io_in_config_0 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_337 = io_in_config_1 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_338 = io_in_config_2 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_339 = io_in_config_3 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_340 = io_in_config_4 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_341 = io_in_config_5 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_342 = io_in_config_6 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_343 = io_in_config_7 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_344 = io_in_config_8 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_345 = io_in_config_9 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_346 = io_in_config_10 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_347 = io_in_config_11 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_348 = io_in_config_12 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_349 = io_in_config_13 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_350 = io_in_config_14 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_351 = io_in_config_15 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_352 = io_in_config_16 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_353 = io_in_config_17 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_354 = io_in_config_18 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_355 = io_in_config_19 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_356 = io_in_config_20 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_357 = io_in_config_21 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_358 = io_in_config_22 == 5'he; // @[FFTDesigns.scala 3194:35]
  wire  _T_360 = io_in_config_0 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_361 = io_in_config_1 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_362 = io_in_config_2 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_363 = io_in_config_3 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_364 = io_in_config_4 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_365 = io_in_config_5 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_366 = io_in_config_6 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_367 = io_in_config_7 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_368 = io_in_config_8 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_369 = io_in_config_9 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_370 = io_in_config_10 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_371 = io_in_config_11 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_372 = io_in_config_12 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_373 = io_in_config_13 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_374 = io_in_config_14 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_375 = io_in_config_15 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_376 = io_in_config_16 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_377 = io_in_config_17 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_378 = io_in_config_18 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_379 = io_in_config_19 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_380 = io_in_config_20 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_381 = io_in_config_21 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_382 = io_in_config_22 == 5'hf; // @[FFTDesigns.scala 3194:35]
  wire  _T_384 = io_in_config_0 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_385 = io_in_config_1 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_386 = io_in_config_2 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_387 = io_in_config_3 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_388 = io_in_config_4 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_389 = io_in_config_5 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_390 = io_in_config_6 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_391 = io_in_config_7 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_392 = io_in_config_8 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_393 = io_in_config_9 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_394 = io_in_config_10 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_395 = io_in_config_11 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_396 = io_in_config_12 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_397 = io_in_config_13 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_398 = io_in_config_14 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_399 = io_in_config_15 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_400 = io_in_config_16 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_401 = io_in_config_17 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_402 = io_in_config_18 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_403 = io_in_config_19 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_404 = io_in_config_20 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_405 = io_in_config_21 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_406 = io_in_config_22 == 5'h10; // @[FFTDesigns.scala 3194:35]
  wire  _T_408 = io_in_config_0 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_409 = io_in_config_1 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_410 = io_in_config_2 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_411 = io_in_config_3 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_412 = io_in_config_4 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_413 = io_in_config_5 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_414 = io_in_config_6 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_415 = io_in_config_7 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_416 = io_in_config_8 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_417 = io_in_config_9 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_418 = io_in_config_10 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_419 = io_in_config_11 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_420 = io_in_config_12 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_421 = io_in_config_13 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_422 = io_in_config_14 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_423 = io_in_config_15 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_424 = io_in_config_16 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_425 = io_in_config_17 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_426 = io_in_config_18 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_427 = io_in_config_19 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_428 = io_in_config_20 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_429 = io_in_config_21 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_430 = io_in_config_22 == 5'h11; // @[FFTDesigns.scala 3194:35]
  wire  _T_432 = io_in_config_0 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_433 = io_in_config_1 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_434 = io_in_config_2 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_435 = io_in_config_3 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_436 = io_in_config_4 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_437 = io_in_config_5 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_438 = io_in_config_6 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_439 = io_in_config_7 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_440 = io_in_config_8 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_441 = io_in_config_9 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_442 = io_in_config_10 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_443 = io_in_config_11 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_444 = io_in_config_12 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_445 = io_in_config_13 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_446 = io_in_config_14 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_447 = io_in_config_15 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_448 = io_in_config_16 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_449 = io_in_config_17 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_450 = io_in_config_18 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_451 = io_in_config_19 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_452 = io_in_config_20 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_453 = io_in_config_21 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_454 = io_in_config_22 == 5'h12; // @[FFTDesigns.scala 3194:35]
  wire  _T_456 = io_in_config_0 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_457 = io_in_config_1 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_458 = io_in_config_2 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_459 = io_in_config_3 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_460 = io_in_config_4 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_461 = io_in_config_5 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_462 = io_in_config_6 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_463 = io_in_config_7 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_464 = io_in_config_8 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_465 = io_in_config_9 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_466 = io_in_config_10 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_467 = io_in_config_11 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_468 = io_in_config_12 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_469 = io_in_config_13 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_470 = io_in_config_14 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_471 = io_in_config_15 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_472 = io_in_config_16 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_473 = io_in_config_17 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_474 = io_in_config_18 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_475 = io_in_config_19 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_476 = io_in_config_20 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_477 = io_in_config_21 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_478 = io_in_config_22 == 5'h13; // @[FFTDesigns.scala 3194:35]
  wire  _T_480 = io_in_config_0 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_481 = io_in_config_1 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_482 = io_in_config_2 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_483 = io_in_config_3 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_484 = io_in_config_4 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_485 = io_in_config_5 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_486 = io_in_config_6 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_487 = io_in_config_7 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_488 = io_in_config_8 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_489 = io_in_config_9 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_490 = io_in_config_10 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_491 = io_in_config_11 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_492 = io_in_config_12 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_493 = io_in_config_13 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_494 = io_in_config_14 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_495 = io_in_config_15 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_496 = io_in_config_16 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_497 = io_in_config_17 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_498 = io_in_config_18 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_499 = io_in_config_19 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_500 = io_in_config_20 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_501 = io_in_config_21 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_502 = io_in_config_22 == 5'h14; // @[FFTDesigns.scala 3194:35]
  wire  _T_504 = io_in_config_0 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_505 = io_in_config_1 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_506 = io_in_config_2 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_507 = io_in_config_3 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_508 = io_in_config_4 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_509 = io_in_config_5 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_510 = io_in_config_6 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_511 = io_in_config_7 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_512 = io_in_config_8 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_513 = io_in_config_9 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_514 = io_in_config_10 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_515 = io_in_config_11 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_516 = io_in_config_12 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_517 = io_in_config_13 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_518 = io_in_config_14 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_519 = io_in_config_15 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_520 = io_in_config_16 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_521 = io_in_config_17 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_522 = io_in_config_18 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_523 = io_in_config_19 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_524 = io_in_config_20 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_525 = io_in_config_21 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_526 = io_in_config_22 == 5'h15; // @[FFTDesigns.scala 3194:35]
  wire  _T_528 = io_in_config_0 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_529 = io_in_config_1 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_530 = io_in_config_2 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_531 = io_in_config_3 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_532 = io_in_config_4 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_533 = io_in_config_5 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_534 = io_in_config_6 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_535 = io_in_config_7 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_536 = io_in_config_8 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_537 = io_in_config_9 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_538 = io_in_config_10 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_539 = io_in_config_11 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_540 = io_in_config_12 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_541 = io_in_config_13 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_542 = io_in_config_14 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_543 = io_in_config_15 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_544 = io_in_config_16 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_545 = io_in_config_17 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_546 = io_in_config_18 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_547 = io_in_config_19 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_548 = io_in_config_20 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_549 = io_in_config_21 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_550 = io_in_config_22 == 5'h16; // @[FFTDesigns.scala 3194:35]
  wire  _T_552 = io_in_config_0 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_553 = io_in_config_1 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_554 = io_in_config_2 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_555 = io_in_config_3 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_556 = io_in_config_4 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_557 = io_in_config_5 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_558 = io_in_config_6 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_559 = io_in_config_7 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_560 = io_in_config_8 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_561 = io_in_config_9 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_562 = io_in_config_10 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_563 = io_in_config_11 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_564 = io_in_config_12 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_565 = io_in_config_13 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_566 = io_in_config_14 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_567 = io_in_config_15 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_568 = io_in_config_16 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_569 = io_in_config_17 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_570 = io_in_config_18 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_571 = io_in_config_19 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_572 = io_in_config_20 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_573 = io_in_config_21 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire  _T_574 = io_in_config_22 == 5'h17; // @[FFTDesigns.scala 3194:35]
  wire [4:0] _pms_pmx_T = _T_22 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_1 = _T_21 ? 5'h15 : _pms_pmx_T; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_2 = _T_20 ? 5'h14 : _pms_pmx_T_1; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_3 = _T_19 ? 5'h13 : _pms_pmx_T_2; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_4 = _T_18 ? 5'h12 : _pms_pmx_T_3; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_5 = _T_17 ? 5'h11 : _pms_pmx_T_4; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_6 = _T_16 ? 5'h10 : _pms_pmx_T_5; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_7 = _T_15 ? 5'hf : _pms_pmx_T_6; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_8 = _T_14 ? 5'he : _pms_pmx_T_7; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_9 = _T_13 ? 5'hd : _pms_pmx_T_8; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_10 = _T_12 ? 5'hc : _pms_pmx_T_9; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_11 = _T_11 ? 5'hb : _pms_pmx_T_10; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_12 = _T_10 ? 5'ha : _pms_pmx_T_11; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_13 = _T_9 ? 5'h9 : _pms_pmx_T_12; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_14 = _T_8 ? 5'h8 : _pms_pmx_T_13; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_15 = _T_7 ? 5'h7 : _pms_pmx_T_14; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_16 = _T_6 ? 5'h6 : _pms_pmx_T_15; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_17 = _T_5 ? 5'h5 : _pms_pmx_T_16; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_18 = _T_4 ? 5'h4 : _pms_pmx_T_17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_19 = _T_3 ? 5'h3 : _pms_pmx_T_18; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_20 = _T_2 ? 5'h2 : _pms_pmx_T_19; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_21 = _T_1 ? 5'h1 : _pms_pmx_T_20; // @[Mux.scala 47:70]
  wire [4:0] pms_0 = _T ? 5'h0 : _pms_pmx_T_21; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_22 = _T_46 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_23 = _T_45 ? 5'h15 : _pms_pmx_T_22; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_24 = _T_44 ? 5'h14 : _pms_pmx_T_23; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_25 = _T_43 ? 5'h13 : _pms_pmx_T_24; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_26 = _T_42 ? 5'h12 : _pms_pmx_T_25; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_27 = _T_41 ? 5'h11 : _pms_pmx_T_26; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_28 = _T_40 ? 5'h10 : _pms_pmx_T_27; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_29 = _T_39 ? 5'hf : _pms_pmx_T_28; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_30 = _T_38 ? 5'he : _pms_pmx_T_29; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_31 = _T_37 ? 5'hd : _pms_pmx_T_30; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_32 = _T_36 ? 5'hc : _pms_pmx_T_31; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_33 = _T_35 ? 5'hb : _pms_pmx_T_32; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_34 = _T_34 ? 5'ha : _pms_pmx_T_33; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_35 = _T_33 ? 5'h9 : _pms_pmx_T_34; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_36 = _T_32 ? 5'h8 : _pms_pmx_T_35; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_37 = _T_31 ? 5'h7 : _pms_pmx_T_36; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_38 = _T_30 ? 5'h6 : _pms_pmx_T_37; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_39 = _T_29 ? 5'h5 : _pms_pmx_T_38; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_40 = _T_28 ? 5'h4 : _pms_pmx_T_39; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_41 = _T_27 ? 5'h3 : _pms_pmx_T_40; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_42 = _T_26 ? 5'h2 : _pms_pmx_T_41; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_43 = _T_25 ? 5'h1 : _pms_pmx_T_42; // @[Mux.scala 47:70]
  wire [4:0] pms_1 = _T_24 ? 5'h0 : _pms_pmx_T_43; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_44 = _T_70 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_45 = _T_69 ? 5'h15 : _pms_pmx_T_44; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_46 = _T_68 ? 5'h14 : _pms_pmx_T_45; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_47 = _T_67 ? 5'h13 : _pms_pmx_T_46; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_48 = _T_66 ? 5'h12 : _pms_pmx_T_47; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_49 = _T_65 ? 5'h11 : _pms_pmx_T_48; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_50 = _T_64 ? 5'h10 : _pms_pmx_T_49; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_51 = _T_63 ? 5'hf : _pms_pmx_T_50; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_52 = _T_62 ? 5'he : _pms_pmx_T_51; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_53 = _T_61 ? 5'hd : _pms_pmx_T_52; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_54 = _T_60 ? 5'hc : _pms_pmx_T_53; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_55 = _T_59 ? 5'hb : _pms_pmx_T_54; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_56 = _T_58 ? 5'ha : _pms_pmx_T_55; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_57 = _T_57 ? 5'h9 : _pms_pmx_T_56; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_58 = _T_56 ? 5'h8 : _pms_pmx_T_57; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_59 = _T_55 ? 5'h7 : _pms_pmx_T_58; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_60 = _T_54 ? 5'h6 : _pms_pmx_T_59; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_61 = _T_53 ? 5'h5 : _pms_pmx_T_60; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_62 = _T_52 ? 5'h4 : _pms_pmx_T_61; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_63 = _T_51 ? 5'h3 : _pms_pmx_T_62; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_64 = _T_50 ? 5'h2 : _pms_pmx_T_63; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_65 = _T_49 ? 5'h1 : _pms_pmx_T_64; // @[Mux.scala 47:70]
  wire [4:0] pms_2 = _T_48 ? 5'h0 : _pms_pmx_T_65; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_66 = _T_94 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_67 = _T_93 ? 5'h15 : _pms_pmx_T_66; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_68 = _T_92 ? 5'h14 : _pms_pmx_T_67; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_69 = _T_91 ? 5'h13 : _pms_pmx_T_68; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_70 = _T_90 ? 5'h12 : _pms_pmx_T_69; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_71 = _T_89 ? 5'h11 : _pms_pmx_T_70; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_72 = _T_88 ? 5'h10 : _pms_pmx_T_71; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_73 = _T_87 ? 5'hf : _pms_pmx_T_72; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_74 = _T_86 ? 5'he : _pms_pmx_T_73; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_75 = _T_85 ? 5'hd : _pms_pmx_T_74; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_76 = _T_84 ? 5'hc : _pms_pmx_T_75; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_77 = _T_83 ? 5'hb : _pms_pmx_T_76; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_78 = _T_82 ? 5'ha : _pms_pmx_T_77; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_79 = _T_81 ? 5'h9 : _pms_pmx_T_78; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_80 = _T_80 ? 5'h8 : _pms_pmx_T_79; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_81 = _T_79 ? 5'h7 : _pms_pmx_T_80; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_82 = _T_78 ? 5'h6 : _pms_pmx_T_81; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_83 = _T_77 ? 5'h5 : _pms_pmx_T_82; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_84 = _T_76 ? 5'h4 : _pms_pmx_T_83; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_85 = _T_75 ? 5'h3 : _pms_pmx_T_84; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_86 = _T_74 ? 5'h2 : _pms_pmx_T_85; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_87 = _T_73 ? 5'h1 : _pms_pmx_T_86; // @[Mux.scala 47:70]
  wire [4:0] pms_3 = _T_72 ? 5'h0 : _pms_pmx_T_87; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_88 = _T_118 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_89 = _T_117 ? 5'h15 : _pms_pmx_T_88; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_90 = _T_116 ? 5'h14 : _pms_pmx_T_89; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_91 = _T_115 ? 5'h13 : _pms_pmx_T_90; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_92 = _T_114 ? 5'h12 : _pms_pmx_T_91; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_93 = _T_113 ? 5'h11 : _pms_pmx_T_92; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_94 = _T_112 ? 5'h10 : _pms_pmx_T_93; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_95 = _T_111 ? 5'hf : _pms_pmx_T_94; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_96 = _T_110 ? 5'he : _pms_pmx_T_95; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_97 = _T_109 ? 5'hd : _pms_pmx_T_96; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_98 = _T_108 ? 5'hc : _pms_pmx_T_97; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_99 = _T_107 ? 5'hb : _pms_pmx_T_98; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_100 = _T_106 ? 5'ha : _pms_pmx_T_99; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_101 = _T_105 ? 5'h9 : _pms_pmx_T_100; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_102 = _T_104 ? 5'h8 : _pms_pmx_T_101; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_103 = _T_103 ? 5'h7 : _pms_pmx_T_102; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_104 = _T_102 ? 5'h6 : _pms_pmx_T_103; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_105 = _T_101 ? 5'h5 : _pms_pmx_T_104; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_106 = _T_100 ? 5'h4 : _pms_pmx_T_105; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_107 = _T_99 ? 5'h3 : _pms_pmx_T_106; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_108 = _T_98 ? 5'h2 : _pms_pmx_T_107; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_109 = _T_97 ? 5'h1 : _pms_pmx_T_108; // @[Mux.scala 47:70]
  wire [4:0] pms_4 = _T_96 ? 5'h0 : _pms_pmx_T_109; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_110 = _T_142 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_111 = _T_141 ? 5'h15 : _pms_pmx_T_110; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_112 = _T_140 ? 5'h14 : _pms_pmx_T_111; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_113 = _T_139 ? 5'h13 : _pms_pmx_T_112; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_114 = _T_138 ? 5'h12 : _pms_pmx_T_113; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_115 = _T_137 ? 5'h11 : _pms_pmx_T_114; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_116 = _T_136 ? 5'h10 : _pms_pmx_T_115; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_117 = _T_135 ? 5'hf : _pms_pmx_T_116; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_118 = _T_134 ? 5'he : _pms_pmx_T_117; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_119 = _T_133 ? 5'hd : _pms_pmx_T_118; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_120 = _T_132 ? 5'hc : _pms_pmx_T_119; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_121 = _T_131 ? 5'hb : _pms_pmx_T_120; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_122 = _T_130 ? 5'ha : _pms_pmx_T_121; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_123 = _T_129 ? 5'h9 : _pms_pmx_T_122; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_124 = _T_128 ? 5'h8 : _pms_pmx_T_123; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_125 = _T_127 ? 5'h7 : _pms_pmx_T_124; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_126 = _T_126 ? 5'h6 : _pms_pmx_T_125; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_127 = _T_125 ? 5'h5 : _pms_pmx_T_126; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_128 = _T_124 ? 5'h4 : _pms_pmx_T_127; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_129 = _T_123 ? 5'h3 : _pms_pmx_T_128; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_130 = _T_122 ? 5'h2 : _pms_pmx_T_129; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_131 = _T_121 ? 5'h1 : _pms_pmx_T_130; // @[Mux.scala 47:70]
  wire [4:0] pms_5 = _T_120 ? 5'h0 : _pms_pmx_T_131; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_132 = _T_166 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_133 = _T_165 ? 5'h15 : _pms_pmx_T_132; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_134 = _T_164 ? 5'h14 : _pms_pmx_T_133; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_135 = _T_163 ? 5'h13 : _pms_pmx_T_134; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_136 = _T_162 ? 5'h12 : _pms_pmx_T_135; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_137 = _T_161 ? 5'h11 : _pms_pmx_T_136; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_138 = _T_160 ? 5'h10 : _pms_pmx_T_137; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_139 = _T_159 ? 5'hf : _pms_pmx_T_138; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_140 = _T_158 ? 5'he : _pms_pmx_T_139; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_141 = _T_157 ? 5'hd : _pms_pmx_T_140; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_142 = _T_156 ? 5'hc : _pms_pmx_T_141; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_143 = _T_155 ? 5'hb : _pms_pmx_T_142; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_144 = _T_154 ? 5'ha : _pms_pmx_T_143; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_145 = _T_153 ? 5'h9 : _pms_pmx_T_144; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_146 = _T_152 ? 5'h8 : _pms_pmx_T_145; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_147 = _T_151 ? 5'h7 : _pms_pmx_T_146; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_148 = _T_150 ? 5'h6 : _pms_pmx_T_147; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_149 = _T_149 ? 5'h5 : _pms_pmx_T_148; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_150 = _T_148 ? 5'h4 : _pms_pmx_T_149; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_151 = _T_147 ? 5'h3 : _pms_pmx_T_150; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_152 = _T_146 ? 5'h2 : _pms_pmx_T_151; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_153 = _T_145 ? 5'h1 : _pms_pmx_T_152; // @[Mux.scala 47:70]
  wire [4:0] pms_6 = _T_144 ? 5'h0 : _pms_pmx_T_153; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_154 = _T_190 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_155 = _T_189 ? 5'h15 : _pms_pmx_T_154; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_156 = _T_188 ? 5'h14 : _pms_pmx_T_155; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_157 = _T_187 ? 5'h13 : _pms_pmx_T_156; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_158 = _T_186 ? 5'h12 : _pms_pmx_T_157; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_159 = _T_185 ? 5'h11 : _pms_pmx_T_158; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_160 = _T_184 ? 5'h10 : _pms_pmx_T_159; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_161 = _T_183 ? 5'hf : _pms_pmx_T_160; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_162 = _T_182 ? 5'he : _pms_pmx_T_161; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_163 = _T_181 ? 5'hd : _pms_pmx_T_162; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_164 = _T_180 ? 5'hc : _pms_pmx_T_163; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_165 = _T_179 ? 5'hb : _pms_pmx_T_164; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_166 = _T_178 ? 5'ha : _pms_pmx_T_165; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_167 = _T_177 ? 5'h9 : _pms_pmx_T_166; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_168 = _T_176 ? 5'h8 : _pms_pmx_T_167; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_169 = _T_175 ? 5'h7 : _pms_pmx_T_168; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_170 = _T_174 ? 5'h6 : _pms_pmx_T_169; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_171 = _T_173 ? 5'h5 : _pms_pmx_T_170; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_172 = _T_172 ? 5'h4 : _pms_pmx_T_171; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_173 = _T_171 ? 5'h3 : _pms_pmx_T_172; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_174 = _T_170 ? 5'h2 : _pms_pmx_T_173; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_175 = _T_169 ? 5'h1 : _pms_pmx_T_174; // @[Mux.scala 47:70]
  wire [4:0] pms_7 = _T_168 ? 5'h0 : _pms_pmx_T_175; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_176 = _T_214 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_177 = _T_213 ? 5'h15 : _pms_pmx_T_176; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_178 = _T_212 ? 5'h14 : _pms_pmx_T_177; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_179 = _T_211 ? 5'h13 : _pms_pmx_T_178; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_180 = _T_210 ? 5'h12 : _pms_pmx_T_179; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_181 = _T_209 ? 5'h11 : _pms_pmx_T_180; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_182 = _T_208 ? 5'h10 : _pms_pmx_T_181; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_183 = _T_207 ? 5'hf : _pms_pmx_T_182; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_184 = _T_206 ? 5'he : _pms_pmx_T_183; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_185 = _T_205 ? 5'hd : _pms_pmx_T_184; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_186 = _T_204 ? 5'hc : _pms_pmx_T_185; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_187 = _T_203 ? 5'hb : _pms_pmx_T_186; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_188 = _T_202 ? 5'ha : _pms_pmx_T_187; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_189 = _T_201 ? 5'h9 : _pms_pmx_T_188; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_190 = _T_200 ? 5'h8 : _pms_pmx_T_189; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_191 = _T_199 ? 5'h7 : _pms_pmx_T_190; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_192 = _T_198 ? 5'h6 : _pms_pmx_T_191; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_193 = _T_197 ? 5'h5 : _pms_pmx_T_192; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_194 = _T_196 ? 5'h4 : _pms_pmx_T_193; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_195 = _T_195 ? 5'h3 : _pms_pmx_T_194; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_196 = _T_194 ? 5'h2 : _pms_pmx_T_195; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_197 = _T_193 ? 5'h1 : _pms_pmx_T_196; // @[Mux.scala 47:70]
  wire [4:0] pms_8 = _T_192 ? 5'h0 : _pms_pmx_T_197; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_198 = _T_238 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_199 = _T_237 ? 5'h15 : _pms_pmx_T_198; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_200 = _T_236 ? 5'h14 : _pms_pmx_T_199; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_201 = _T_235 ? 5'h13 : _pms_pmx_T_200; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_202 = _T_234 ? 5'h12 : _pms_pmx_T_201; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_203 = _T_233 ? 5'h11 : _pms_pmx_T_202; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_204 = _T_232 ? 5'h10 : _pms_pmx_T_203; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_205 = _T_231 ? 5'hf : _pms_pmx_T_204; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_206 = _T_230 ? 5'he : _pms_pmx_T_205; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_207 = _T_229 ? 5'hd : _pms_pmx_T_206; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_208 = _T_228 ? 5'hc : _pms_pmx_T_207; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_209 = _T_227 ? 5'hb : _pms_pmx_T_208; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_210 = _T_226 ? 5'ha : _pms_pmx_T_209; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_211 = _T_225 ? 5'h9 : _pms_pmx_T_210; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_212 = _T_224 ? 5'h8 : _pms_pmx_T_211; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_213 = _T_223 ? 5'h7 : _pms_pmx_T_212; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_214 = _T_222 ? 5'h6 : _pms_pmx_T_213; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_215 = _T_221 ? 5'h5 : _pms_pmx_T_214; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_216 = _T_220 ? 5'h4 : _pms_pmx_T_215; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_217 = _T_219 ? 5'h3 : _pms_pmx_T_216; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_218 = _T_218 ? 5'h2 : _pms_pmx_T_217; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_219 = _T_217 ? 5'h1 : _pms_pmx_T_218; // @[Mux.scala 47:70]
  wire [4:0] pms_9 = _T_216 ? 5'h0 : _pms_pmx_T_219; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_220 = _T_262 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_221 = _T_261 ? 5'h15 : _pms_pmx_T_220; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_222 = _T_260 ? 5'h14 : _pms_pmx_T_221; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_223 = _T_259 ? 5'h13 : _pms_pmx_T_222; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_224 = _T_258 ? 5'h12 : _pms_pmx_T_223; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_225 = _T_257 ? 5'h11 : _pms_pmx_T_224; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_226 = _T_256 ? 5'h10 : _pms_pmx_T_225; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_227 = _T_255 ? 5'hf : _pms_pmx_T_226; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_228 = _T_254 ? 5'he : _pms_pmx_T_227; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_229 = _T_253 ? 5'hd : _pms_pmx_T_228; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_230 = _T_252 ? 5'hc : _pms_pmx_T_229; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_231 = _T_251 ? 5'hb : _pms_pmx_T_230; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_232 = _T_250 ? 5'ha : _pms_pmx_T_231; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_233 = _T_249 ? 5'h9 : _pms_pmx_T_232; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_234 = _T_248 ? 5'h8 : _pms_pmx_T_233; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_235 = _T_247 ? 5'h7 : _pms_pmx_T_234; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_236 = _T_246 ? 5'h6 : _pms_pmx_T_235; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_237 = _T_245 ? 5'h5 : _pms_pmx_T_236; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_238 = _T_244 ? 5'h4 : _pms_pmx_T_237; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_239 = _T_243 ? 5'h3 : _pms_pmx_T_238; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_240 = _T_242 ? 5'h2 : _pms_pmx_T_239; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_241 = _T_241 ? 5'h1 : _pms_pmx_T_240; // @[Mux.scala 47:70]
  wire [4:0] pms_10 = _T_240 ? 5'h0 : _pms_pmx_T_241; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_242 = _T_286 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_243 = _T_285 ? 5'h15 : _pms_pmx_T_242; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_244 = _T_284 ? 5'h14 : _pms_pmx_T_243; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_245 = _T_283 ? 5'h13 : _pms_pmx_T_244; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_246 = _T_282 ? 5'h12 : _pms_pmx_T_245; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_247 = _T_281 ? 5'h11 : _pms_pmx_T_246; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_248 = _T_280 ? 5'h10 : _pms_pmx_T_247; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_249 = _T_279 ? 5'hf : _pms_pmx_T_248; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_250 = _T_278 ? 5'he : _pms_pmx_T_249; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_251 = _T_277 ? 5'hd : _pms_pmx_T_250; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_252 = _T_276 ? 5'hc : _pms_pmx_T_251; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_253 = _T_275 ? 5'hb : _pms_pmx_T_252; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_254 = _T_274 ? 5'ha : _pms_pmx_T_253; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_255 = _T_273 ? 5'h9 : _pms_pmx_T_254; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_256 = _T_272 ? 5'h8 : _pms_pmx_T_255; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_257 = _T_271 ? 5'h7 : _pms_pmx_T_256; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_258 = _T_270 ? 5'h6 : _pms_pmx_T_257; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_259 = _T_269 ? 5'h5 : _pms_pmx_T_258; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_260 = _T_268 ? 5'h4 : _pms_pmx_T_259; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_261 = _T_267 ? 5'h3 : _pms_pmx_T_260; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_262 = _T_266 ? 5'h2 : _pms_pmx_T_261; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_263 = _T_265 ? 5'h1 : _pms_pmx_T_262; // @[Mux.scala 47:70]
  wire [4:0] pms_11 = _T_264 ? 5'h0 : _pms_pmx_T_263; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_264 = _T_310 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_265 = _T_309 ? 5'h15 : _pms_pmx_T_264; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_266 = _T_308 ? 5'h14 : _pms_pmx_T_265; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_267 = _T_307 ? 5'h13 : _pms_pmx_T_266; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_268 = _T_306 ? 5'h12 : _pms_pmx_T_267; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_269 = _T_305 ? 5'h11 : _pms_pmx_T_268; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_270 = _T_304 ? 5'h10 : _pms_pmx_T_269; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_271 = _T_303 ? 5'hf : _pms_pmx_T_270; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_272 = _T_302 ? 5'he : _pms_pmx_T_271; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_273 = _T_301 ? 5'hd : _pms_pmx_T_272; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_274 = _T_300 ? 5'hc : _pms_pmx_T_273; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_275 = _T_299 ? 5'hb : _pms_pmx_T_274; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_276 = _T_298 ? 5'ha : _pms_pmx_T_275; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_277 = _T_297 ? 5'h9 : _pms_pmx_T_276; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_278 = _T_296 ? 5'h8 : _pms_pmx_T_277; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_279 = _T_295 ? 5'h7 : _pms_pmx_T_278; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_280 = _T_294 ? 5'h6 : _pms_pmx_T_279; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_281 = _T_293 ? 5'h5 : _pms_pmx_T_280; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_282 = _T_292 ? 5'h4 : _pms_pmx_T_281; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_283 = _T_291 ? 5'h3 : _pms_pmx_T_282; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_284 = _T_290 ? 5'h2 : _pms_pmx_T_283; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_285 = _T_289 ? 5'h1 : _pms_pmx_T_284; // @[Mux.scala 47:70]
  wire [4:0] pms_12 = _T_288 ? 5'h0 : _pms_pmx_T_285; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_286 = _T_334 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_287 = _T_333 ? 5'h15 : _pms_pmx_T_286; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_288 = _T_332 ? 5'h14 : _pms_pmx_T_287; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_289 = _T_331 ? 5'h13 : _pms_pmx_T_288; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_290 = _T_330 ? 5'h12 : _pms_pmx_T_289; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_291 = _T_329 ? 5'h11 : _pms_pmx_T_290; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_292 = _T_328 ? 5'h10 : _pms_pmx_T_291; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_293 = _T_327 ? 5'hf : _pms_pmx_T_292; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_294 = _T_326 ? 5'he : _pms_pmx_T_293; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_295 = _T_325 ? 5'hd : _pms_pmx_T_294; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_296 = _T_324 ? 5'hc : _pms_pmx_T_295; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_297 = _T_323 ? 5'hb : _pms_pmx_T_296; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_298 = _T_322 ? 5'ha : _pms_pmx_T_297; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_299 = _T_321 ? 5'h9 : _pms_pmx_T_298; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_300 = _T_320 ? 5'h8 : _pms_pmx_T_299; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_301 = _T_319 ? 5'h7 : _pms_pmx_T_300; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_302 = _T_318 ? 5'h6 : _pms_pmx_T_301; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_303 = _T_317 ? 5'h5 : _pms_pmx_T_302; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_304 = _T_316 ? 5'h4 : _pms_pmx_T_303; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_305 = _T_315 ? 5'h3 : _pms_pmx_T_304; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_306 = _T_314 ? 5'h2 : _pms_pmx_T_305; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_307 = _T_313 ? 5'h1 : _pms_pmx_T_306; // @[Mux.scala 47:70]
  wire [4:0] pms_13 = _T_312 ? 5'h0 : _pms_pmx_T_307; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_308 = _T_358 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_309 = _T_357 ? 5'h15 : _pms_pmx_T_308; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_310 = _T_356 ? 5'h14 : _pms_pmx_T_309; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_311 = _T_355 ? 5'h13 : _pms_pmx_T_310; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_312 = _T_354 ? 5'h12 : _pms_pmx_T_311; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_313 = _T_353 ? 5'h11 : _pms_pmx_T_312; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_314 = _T_352 ? 5'h10 : _pms_pmx_T_313; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_315 = _T_351 ? 5'hf : _pms_pmx_T_314; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_316 = _T_350 ? 5'he : _pms_pmx_T_315; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_317 = _T_349 ? 5'hd : _pms_pmx_T_316; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_318 = _T_348 ? 5'hc : _pms_pmx_T_317; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_319 = _T_347 ? 5'hb : _pms_pmx_T_318; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_320 = _T_346 ? 5'ha : _pms_pmx_T_319; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_321 = _T_345 ? 5'h9 : _pms_pmx_T_320; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_322 = _T_344 ? 5'h8 : _pms_pmx_T_321; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_323 = _T_343 ? 5'h7 : _pms_pmx_T_322; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_324 = _T_342 ? 5'h6 : _pms_pmx_T_323; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_325 = _T_341 ? 5'h5 : _pms_pmx_T_324; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_326 = _T_340 ? 5'h4 : _pms_pmx_T_325; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_327 = _T_339 ? 5'h3 : _pms_pmx_T_326; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_328 = _T_338 ? 5'h2 : _pms_pmx_T_327; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_329 = _T_337 ? 5'h1 : _pms_pmx_T_328; // @[Mux.scala 47:70]
  wire [4:0] pms_14 = _T_336 ? 5'h0 : _pms_pmx_T_329; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_330 = _T_382 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_331 = _T_381 ? 5'h15 : _pms_pmx_T_330; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_332 = _T_380 ? 5'h14 : _pms_pmx_T_331; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_333 = _T_379 ? 5'h13 : _pms_pmx_T_332; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_334 = _T_378 ? 5'h12 : _pms_pmx_T_333; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_335 = _T_377 ? 5'h11 : _pms_pmx_T_334; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_336 = _T_376 ? 5'h10 : _pms_pmx_T_335; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_337 = _T_375 ? 5'hf : _pms_pmx_T_336; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_338 = _T_374 ? 5'he : _pms_pmx_T_337; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_339 = _T_373 ? 5'hd : _pms_pmx_T_338; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_340 = _T_372 ? 5'hc : _pms_pmx_T_339; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_341 = _T_371 ? 5'hb : _pms_pmx_T_340; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_342 = _T_370 ? 5'ha : _pms_pmx_T_341; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_343 = _T_369 ? 5'h9 : _pms_pmx_T_342; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_344 = _T_368 ? 5'h8 : _pms_pmx_T_343; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_345 = _T_367 ? 5'h7 : _pms_pmx_T_344; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_346 = _T_366 ? 5'h6 : _pms_pmx_T_345; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_347 = _T_365 ? 5'h5 : _pms_pmx_T_346; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_348 = _T_364 ? 5'h4 : _pms_pmx_T_347; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_349 = _T_363 ? 5'h3 : _pms_pmx_T_348; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_350 = _T_362 ? 5'h2 : _pms_pmx_T_349; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_351 = _T_361 ? 5'h1 : _pms_pmx_T_350; // @[Mux.scala 47:70]
  wire [4:0] pms_15 = _T_360 ? 5'h0 : _pms_pmx_T_351; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_352 = _T_406 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_353 = _T_405 ? 5'h15 : _pms_pmx_T_352; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_354 = _T_404 ? 5'h14 : _pms_pmx_T_353; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_355 = _T_403 ? 5'h13 : _pms_pmx_T_354; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_356 = _T_402 ? 5'h12 : _pms_pmx_T_355; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_357 = _T_401 ? 5'h11 : _pms_pmx_T_356; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_358 = _T_400 ? 5'h10 : _pms_pmx_T_357; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_359 = _T_399 ? 5'hf : _pms_pmx_T_358; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_360 = _T_398 ? 5'he : _pms_pmx_T_359; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_361 = _T_397 ? 5'hd : _pms_pmx_T_360; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_362 = _T_396 ? 5'hc : _pms_pmx_T_361; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_363 = _T_395 ? 5'hb : _pms_pmx_T_362; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_364 = _T_394 ? 5'ha : _pms_pmx_T_363; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_365 = _T_393 ? 5'h9 : _pms_pmx_T_364; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_366 = _T_392 ? 5'h8 : _pms_pmx_T_365; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_367 = _T_391 ? 5'h7 : _pms_pmx_T_366; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_368 = _T_390 ? 5'h6 : _pms_pmx_T_367; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_369 = _T_389 ? 5'h5 : _pms_pmx_T_368; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_370 = _T_388 ? 5'h4 : _pms_pmx_T_369; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_371 = _T_387 ? 5'h3 : _pms_pmx_T_370; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_372 = _T_386 ? 5'h2 : _pms_pmx_T_371; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_373 = _T_385 ? 5'h1 : _pms_pmx_T_372; // @[Mux.scala 47:70]
  wire [4:0] pms_16 = _T_384 ? 5'h0 : _pms_pmx_T_373; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_374 = _T_430 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_375 = _T_429 ? 5'h15 : _pms_pmx_T_374; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_376 = _T_428 ? 5'h14 : _pms_pmx_T_375; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_377 = _T_427 ? 5'h13 : _pms_pmx_T_376; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_378 = _T_426 ? 5'h12 : _pms_pmx_T_377; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_379 = _T_425 ? 5'h11 : _pms_pmx_T_378; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_380 = _T_424 ? 5'h10 : _pms_pmx_T_379; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_381 = _T_423 ? 5'hf : _pms_pmx_T_380; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_382 = _T_422 ? 5'he : _pms_pmx_T_381; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_383 = _T_421 ? 5'hd : _pms_pmx_T_382; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_384 = _T_420 ? 5'hc : _pms_pmx_T_383; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_385 = _T_419 ? 5'hb : _pms_pmx_T_384; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_386 = _T_418 ? 5'ha : _pms_pmx_T_385; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_387 = _T_417 ? 5'h9 : _pms_pmx_T_386; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_388 = _T_416 ? 5'h8 : _pms_pmx_T_387; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_389 = _T_415 ? 5'h7 : _pms_pmx_T_388; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_390 = _T_414 ? 5'h6 : _pms_pmx_T_389; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_391 = _T_413 ? 5'h5 : _pms_pmx_T_390; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_392 = _T_412 ? 5'h4 : _pms_pmx_T_391; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_393 = _T_411 ? 5'h3 : _pms_pmx_T_392; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_394 = _T_410 ? 5'h2 : _pms_pmx_T_393; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_395 = _T_409 ? 5'h1 : _pms_pmx_T_394; // @[Mux.scala 47:70]
  wire [4:0] pms_17 = _T_408 ? 5'h0 : _pms_pmx_T_395; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_396 = _T_454 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_397 = _T_453 ? 5'h15 : _pms_pmx_T_396; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_398 = _T_452 ? 5'h14 : _pms_pmx_T_397; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_399 = _T_451 ? 5'h13 : _pms_pmx_T_398; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_400 = _T_450 ? 5'h12 : _pms_pmx_T_399; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_401 = _T_449 ? 5'h11 : _pms_pmx_T_400; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_402 = _T_448 ? 5'h10 : _pms_pmx_T_401; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_403 = _T_447 ? 5'hf : _pms_pmx_T_402; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_404 = _T_446 ? 5'he : _pms_pmx_T_403; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_405 = _T_445 ? 5'hd : _pms_pmx_T_404; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_406 = _T_444 ? 5'hc : _pms_pmx_T_405; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_407 = _T_443 ? 5'hb : _pms_pmx_T_406; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_408 = _T_442 ? 5'ha : _pms_pmx_T_407; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_409 = _T_441 ? 5'h9 : _pms_pmx_T_408; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_410 = _T_440 ? 5'h8 : _pms_pmx_T_409; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_411 = _T_439 ? 5'h7 : _pms_pmx_T_410; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_412 = _T_438 ? 5'h6 : _pms_pmx_T_411; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_413 = _T_437 ? 5'h5 : _pms_pmx_T_412; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_414 = _T_436 ? 5'h4 : _pms_pmx_T_413; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_415 = _T_435 ? 5'h3 : _pms_pmx_T_414; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_416 = _T_434 ? 5'h2 : _pms_pmx_T_415; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_417 = _T_433 ? 5'h1 : _pms_pmx_T_416; // @[Mux.scala 47:70]
  wire [4:0] pms_18 = _T_432 ? 5'h0 : _pms_pmx_T_417; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_418 = _T_478 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_419 = _T_477 ? 5'h15 : _pms_pmx_T_418; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_420 = _T_476 ? 5'h14 : _pms_pmx_T_419; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_421 = _T_475 ? 5'h13 : _pms_pmx_T_420; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_422 = _T_474 ? 5'h12 : _pms_pmx_T_421; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_423 = _T_473 ? 5'h11 : _pms_pmx_T_422; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_424 = _T_472 ? 5'h10 : _pms_pmx_T_423; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_425 = _T_471 ? 5'hf : _pms_pmx_T_424; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_426 = _T_470 ? 5'he : _pms_pmx_T_425; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_427 = _T_469 ? 5'hd : _pms_pmx_T_426; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_428 = _T_468 ? 5'hc : _pms_pmx_T_427; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_429 = _T_467 ? 5'hb : _pms_pmx_T_428; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_430 = _T_466 ? 5'ha : _pms_pmx_T_429; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_431 = _T_465 ? 5'h9 : _pms_pmx_T_430; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_432 = _T_464 ? 5'h8 : _pms_pmx_T_431; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_433 = _T_463 ? 5'h7 : _pms_pmx_T_432; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_434 = _T_462 ? 5'h6 : _pms_pmx_T_433; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_435 = _T_461 ? 5'h5 : _pms_pmx_T_434; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_436 = _T_460 ? 5'h4 : _pms_pmx_T_435; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_437 = _T_459 ? 5'h3 : _pms_pmx_T_436; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_438 = _T_458 ? 5'h2 : _pms_pmx_T_437; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_439 = _T_457 ? 5'h1 : _pms_pmx_T_438; // @[Mux.scala 47:70]
  wire [4:0] pms_19 = _T_456 ? 5'h0 : _pms_pmx_T_439; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_440 = _T_502 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_441 = _T_501 ? 5'h15 : _pms_pmx_T_440; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_442 = _T_500 ? 5'h14 : _pms_pmx_T_441; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_443 = _T_499 ? 5'h13 : _pms_pmx_T_442; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_444 = _T_498 ? 5'h12 : _pms_pmx_T_443; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_445 = _T_497 ? 5'h11 : _pms_pmx_T_444; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_446 = _T_496 ? 5'h10 : _pms_pmx_T_445; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_447 = _T_495 ? 5'hf : _pms_pmx_T_446; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_448 = _T_494 ? 5'he : _pms_pmx_T_447; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_449 = _T_493 ? 5'hd : _pms_pmx_T_448; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_450 = _T_492 ? 5'hc : _pms_pmx_T_449; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_451 = _T_491 ? 5'hb : _pms_pmx_T_450; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_452 = _T_490 ? 5'ha : _pms_pmx_T_451; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_453 = _T_489 ? 5'h9 : _pms_pmx_T_452; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_454 = _T_488 ? 5'h8 : _pms_pmx_T_453; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_455 = _T_487 ? 5'h7 : _pms_pmx_T_454; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_456 = _T_486 ? 5'h6 : _pms_pmx_T_455; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_457 = _T_485 ? 5'h5 : _pms_pmx_T_456; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_458 = _T_484 ? 5'h4 : _pms_pmx_T_457; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_459 = _T_483 ? 5'h3 : _pms_pmx_T_458; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_460 = _T_482 ? 5'h2 : _pms_pmx_T_459; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_461 = _T_481 ? 5'h1 : _pms_pmx_T_460; // @[Mux.scala 47:70]
  wire [4:0] pms_20 = _T_480 ? 5'h0 : _pms_pmx_T_461; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_462 = _T_526 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_463 = _T_525 ? 5'h15 : _pms_pmx_T_462; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_464 = _T_524 ? 5'h14 : _pms_pmx_T_463; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_465 = _T_523 ? 5'h13 : _pms_pmx_T_464; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_466 = _T_522 ? 5'h12 : _pms_pmx_T_465; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_467 = _T_521 ? 5'h11 : _pms_pmx_T_466; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_468 = _T_520 ? 5'h10 : _pms_pmx_T_467; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_469 = _T_519 ? 5'hf : _pms_pmx_T_468; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_470 = _T_518 ? 5'he : _pms_pmx_T_469; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_471 = _T_517 ? 5'hd : _pms_pmx_T_470; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_472 = _T_516 ? 5'hc : _pms_pmx_T_471; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_473 = _T_515 ? 5'hb : _pms_pmx_T_472; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_474 = _T_514 ? 5'ha : _pms_pmx_T_473; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_475 = _T_513 ? 5'h9 : _pms_pmx_T_474; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_476 = _T_512 ? 5'h8 : _pms_pmx_T_475; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_477 = _T_511 ? 5'h7 : _pms_pmx_T_476; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_478 = _T_510 ? 5'h6 : _pms_pmx_T_477; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_479 = _T_509 ? 5'h5 : _pms_pmx_T_478; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_480 = _T_508 ? 5'h4 : _pms_pmx_T_479; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_481 = _T_507 ? 5'h3 : _pms_pmx_T_480; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_482 = _T_506 ? 5'h2 : _pms_pmx_T_481; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_483 = _T_505 ? 5'h1 : _pms_pmx_T_482; // @[Mux.scala 47:70]
  wire [4:0] pms_21 = _T_504 ? 5'h0 : _pms_pmx_T_483; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_484 = _T_550 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_485 = _T_549 ? 5'h15 : _pms_pmx_T_484; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_486 = _T_548 ? 5'h14 : _pms_pmx_T_485; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_487 = _T_547 ? 5'h13 : _pms_pmx_T_486; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_488 = _T_546 ? 5'h12 : _pms_pmx_T_487; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_489 = _T_545 ? 5'h11 : _pms_pmx_T_488; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_490 = _T_544 ? 5'h10 : _pms_pmx_T_489; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_491 = _T_543 ? 5'hf : _pms_pmx_T_490; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_492 = _T_542 ? 5'he : _pms_pmx_T_491; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_493 = _T_541 ? 5'hd : _pms_pmx_T_492; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_494 = _T_540 ? 5'hc : _pms_pmx_T_493; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_495 = _T_539 ? 5'hb : _pms_pmx_T_494; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_496 = _T_538 ? 5'ha : _pms_pmx_T_495; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_497 = _T_537 ? 5'h9 : _pms_pmx_T_496; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_498 = _T_536 ? 5'h8 : _pms_pmx_T_497; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_499 = _T_535 ? 5'h7 : _pms_pmx_T_498; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_500 = _T_534 ? 5'h6 : _pms_pmx_T_499; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_501 = _T_533 ? 5'h5 : _pms_pmx_T_500; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_502 = _T_532 ? 5'h4 : _pms_pmx_T_501; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_503 = _T_531 ? 5'h3 : _pms_pmx_T_502; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_504 = _T_530 ? 5'h2 : _pms_pmx_T_503; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_505 = _T_529 ? 5'h1 : _pms_pmx_T_504; // @[Mux.scala 47:70]
  wire [4:0] pms_22 = _T_528 ? 5'h0 : _pms_pmx_T_505; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_506 = _T_574 ? 5'h16 : 5'h17; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_507 = _T_573 ? 5'h15 : _pms_pmx_T_506; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_508 = _T_572 ? 5'h14 : _pms_pmx_T_507; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_509 = _T_571 ? 5'h13 : _pms_pmx_T_508; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_510 = _T_570 ? 5'h12 : _pms_pmx_T_509; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_511 = _T_569 ? 5'h11 : _pms_pmx_T_510; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_512 = _T_568 ? 5'h10 : _pms_pmx_T_511; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_513 = _T_567 ? 5'hf : _pms_pmx_T_512; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_514 = _T_566 ? 5'he : _pms_pmx_T_513; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_515 = _T_565 ? 5'hd : _pms_pmx_T_514; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_516 = _T_564 ? 5'hc : _pms_pmx_T_515; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_517 = _T_563 ? 5'hb : _pms_pmx_T_516; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_518 = _T_562 ? 5'ha : _pms_pmx_T_517; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_519 = _T_561 ? 5'h9 : _pms_pmx_T_518; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_520 = _T_560 ? 5'h8 : _pms_pmx_T_519; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_521 = _T_559 ? 5'h7 : _pms_pmx_T_520; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_522 = _T_558 ? 5'h6 : _pms_pmx_T_521; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_523 = _T_557 ? 5'h5 : _pms_pmx_T_522; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_524 = _T_556 ? 5'h4 : _pms_pmx_T_523; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_525 = _T_555 ? 5'h3 : _pms_pmx_T_524; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_526 = _T_554 ? 5'h2 : _pms_pmx_T_525; // @[Mux.scala 47:70]
  wire [4:0] _pms_pmx_T_527 = _T_553 ? 5'h1 : _pms_pmx_T_526; // @[Mux.scala 47:70]
  wire [4:0] pms_23 = _T_552 ? 5'h0 : _pms_pmx_T_527; // @[Mux.scala 47:70]
  wire [31:0] _GEN_1 = 5'h1 == pms_0 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_2 = 5'h2 == pms_0 ? io_in_2_Im : _GEN_1; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_3 = 5'h3 == pms_0 ? io_in_3_Im : _GEN_2; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_4 = 5'h4 == pms_0 ? io_in_4_Im : _GEN_3; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_5 = 5'h5 == pms_0 ? io_in_5_Im : _GEN_4; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_6 = 5'h6 == pms_0 ? io_in_6_Im : _GEN_5; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_7 = 5'h7 == pms_0 ? io_in_7_Im : _GEN_6; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_8 = 5'h8 == pms_0 ? io_in_8_Im : _GEN_7; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_9 = 5'h9 == pms_0 ? io_in_9_Im : _GEN_8; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_10 = 5'ha == pms_0 ? io_in_10_Im : _GEN_9; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_11 = 5'hb == pms_0 ? io_in_11_Im : _GEN_10; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_12 = 5'hc == pms_0 ? io_in_12_Im : _GEN_11; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_13 = 5'hd == pms_0 ? io_in_13_Im : _GEN_12; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_14 = 5'he == pms_0 ? io_in_14_Im : _GEN_13; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_15 = 5'hf == pms_0 ? io_in_15_Im : _GEN_14; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_16 = 5'h10 == pms_0 ? io_in_16_Im : _GEN_15; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_17 = 5'h11 == pms_0 ? io_in_17_Im : _GEN_16; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_18 = 5'h12 == pms_0 ? io_in_18_Im : _GEN_17; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_19 = 5'h13 == pms_0 ? io_in_19_Im : _GEN_18; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_20 = 5'h14 == pms_0 ? io_in_20_Im : _GEN_19; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_21 = 5'h15 == pms_0 ? io_in_21_Im : _GEN_20; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_22 = 5'h16 == pms_0 ? io_in_22_Im : _GEN_21; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_25 = 5'h1 == pms_0 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_26 = 5'h2 == pms_0 ? io_in_2_Re : _GEN_25; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_27 = 5'h3 == pms_0 ? io_in_3_Re : _GEN_26; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_28 = 5'h4 == pms_0 ? io_in_4_Re : _GEN_27; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_29 = 5'h5 == pms_0 ? io_in_5_Re : _GEN_28; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_30 = 5'h6 == pms_0 ? io_in_6_Re : _GEN_29; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_31 = 5'h7 == pms_0 ? io_in_7_Re : _GEN_30; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_32 = 5'h8 == pms_0 ? io_in_8_Re : _GEN_31; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_33 = 5'h9 == pms_0 ? io_in_9_Re : _GEN_32; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_34 = 5'ha == pms_0 ? io_in_10_Re : _GEN_33; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_35 = 5'hb == pms_0 ? io_in_11_Re : _GEN_34; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_36 = 5'hc == pms_0 ? io_in_12_Re : _GEN_35; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_37 = 5'hd == pms_0 ? io_in_13_Re : _GEN_36; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_38 = 5'he == pms_0 ? io_in_14_Re : _GEN_37; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_39 = 5'hf == pms_0 ? io_in_15_Re : _GEN_38; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_40 = 5'h10 == pms_0 ? io_in_16_Re : _GEN_39; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_41 = 5'h11 == pms_0 ? io_in_17_Re : _GEN_40; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_42 = 5'h12 == pms_0 ? io_in_18_Re : _GEN_41; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_43 = 5'h13 == pms_0 ? io_in_19_Re : _GEN_42; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_44 = 5'h14 == pms_0 ? io_in_20_Re : _GEN_43; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_45 = 5'h15 == pms_0 ? io_in_21_Re : _GEN_44; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_46 = 5'h16 == pms_0 ? io_in_22_Re : _GEN_45; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_49 = 5'h1 == pms_1 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_50 = 5'h2 == pms_1 ? io_in_2_Im : _GEN_49; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_51 = 5'h3 == pms_1 ? io_in_3_Im : _GEN_50; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_52 = 5'h4 == pms_1 ? io_in_4_Im : _GEN_51; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_53 = 5'h5 == pms_1 ? io_in_5_Im : _GEN_52; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_54 = 5'h6 == pms_1 ? io_in_6_Im : _GEN_53; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_55 = 5'h7 == pms_1 ? io_in_7_Im : _GEN_54; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_56 = 5'h8 == pms_1 ? io_in_8_Im : _GEN_55; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_57 = 5'h9 == pms_1 ? io_in_9_Im : _GEN_56; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_58 = 5'ha == pms_1 ? io_in_10_Im : _GEN_57; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_59 = 5'hb == pms_1 ? io_in_11_Im : _GEN_58; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_60 = 5'hc == pms_1 ? io_in_12_Im : _GEN_59; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_61 = 5'hd == pms_1 ? io_in_13_Im : _GEN_60; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_62 = 5'he == pms_1 ? io_in_14_Im : _GEN_61; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_63 = 5'hf == pms_1 ? io_in_15_Im : _GEN_62; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_64 = 5'h10 == pms_1 ? io_in_16_Im : _GEN_63; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_65 = 5'h11 == pms_1 ? io_in_17_Im : _GEN_64; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_66 = 5'h12 == pms_1 ? io_in_18_Im : _GEN_65; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_67 = 5'h13 == pms_1 ? io_in_19_Im : _GEN_66; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_68 = 5'h14 == pms_1 ? io_in_20_Im : _GEN_67; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_69 = 5'h15 == pms_1 ? io_in_21_Im : _GEN_68; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_70 = 5'h16 == pms_1 ? io_in_22_Im : _GEN_69; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_73 = 5'h1 == pms_1 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_74 = 5'h2 == pms_1 ? io_in_2_Re : _GEN_73; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_75 = 5'h3 == pms_1 ? io_in_3_Re : _GEN_74; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_76 = 5'h4 == pms_1 ? io_in_4_Re : _GEN_75; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_77 = 5'h5 == pms_1 ? io_in_5_Re : _GEN_76; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_78 = 5'h6 == pms_1 ? io_in_6_Re : _GEN_77; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_79 = 5'h7 == pms_1 ? io_in_7_Re : _GEN_78; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_80 = 5'h8 == pms_1 ? io_in_8_Re : _GEN_79; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_81 = 5'h9 == pms_1 ? io_in_9_Re : _GEN_80; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_82 = 5'ha == pms_1 ? io_in_10_Re : _GEN_81; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_83 = 5'hb == pms_1 ? io_in_11_Re : _GEN_82; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_84 = 5'hc == pms_1 ? io_in_12_Re : _GEN_83; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_85 = 5'hd == pms_1 ? io_in_13_Re : _GEN_84; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_86 = 5'he == pms_1 ? io_in_14_Re : _GEN_85; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_87 = 5'hf == pms_1 ? io_in_15_Re : _GEN_86; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_88 = 5'h10 == pms_1 ? io_in_16_Re : _GEN_87; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_89 = 5'h11 == pms_1 ? io_in_17_Re : _GEN_88; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_90 = 5'h12 == pms_1 ? io_in_18_Re : _GEN_89; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_91 = 5'h13 == pms_1 ? io_in_19_Re : _GEN_90; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_92 = 5'h14 == pms_1 ? io_in_20_Re : _GEN_91; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_93 = 5'h15 == pms_1 ? io_in_21_Re : _GEN_92; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_94 = 5'h16 == pms_1 ? io_in_22_Re : _GEN_93; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_97 = 5'h1 == pms_2 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_98 = 5'h2 == pms_2 ? io_in_2_Im : _GEN_97; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_99 = 5'h3 == pms_2 ? io_in_3_Im : _GEN_98; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_100 = 5'h4 == pms_2 ? io_in_4_Im : _GEN_99; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_101 = 5'h5 == pms_2 ? io_in_5_Im : _GEN_100; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_102 = 5'h6 == pms_2 ? io_in_6_Im : _GEN_101; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_103 = 5'h7 == pms_2 ? io_in_7_Im : _GEN_102; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_104 = 5'h8 == pms_2 ? io_in_8_Im : _GEN_103; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_105 = 5'h9 == pms_2 ? io_in_9_Im : _GEN_104; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_106 = 5'ha == pms_2 ? io_in_10_Im : _GEN_105; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_107 = 5'hb == pms_2 ? io_in_11_Im : _GEN_106; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_108 = 5'hc == pms_2 ? io_in_12_Im : _GEN_107; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_109 = 5'hd == pms_2 ? io_in_13_Im : _GEN_108; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_110 = 5'he == pms_2 ? io_in_14_Im : _GEN_109; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_111 = 5'hf == pms_2 ? io_in_15_Im : _GEN_110; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_112 = 5'h10 == pms_2 ? io_in_16_Im : _GEN_111; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_113 = 5'h11 == pms_2 ? io_in_17_Im : _GEN_112; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_114 = 5'h12 == pms_2 ? io_in_18_Im : _GEN_113; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_115 = 5'h13 == pms_2 ? io_in_19_Im : _GEN_114; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_116 = 5'h14 == pms_2 ? io_in_20_Im : _GEN_115; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_117 = 5'h15 == pms_2 ? io_in_21_Im : _GEN_116; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_118 = 5'h16 == pms_2 ? io_in_22_Im : _GEN_117; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_121 = 5'h1 == pms_2 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_122 = 5'h2 == pms_2 ? io_in_2_Re : _GEN_121; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_123 = 5'h3 == pms_2 ? io_in_3_Re : _GEN_122; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_124 = 5'h4 == pms_2 ? io_in_4_Re : _GEN_123; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_125 = 5'h5 == pms_2 ? io_in_5_Re : _GEN_124; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_126 = 5'h6 == pms_2 ? io_in_6_Re : _GEN_125; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_127 = 5'h7 == pms_2 ? io_in_7_Re : _GEN_126; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_128 = 5'h8 == pms_2 ? io_in_8_Re : _GEN_127; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_129 = 5'h9 == pms_2 ? io_in_9_Re : _GEN_128; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_130 = 5'ha == pms_2 ? io_in_10_Re : _GEN_129; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_131 = 5'hb == pms_2 ? io_in_11_Re : _GEN_130; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_132 = 5'hc == pms_2 ? io_in_12_Re : _GEN_131; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_133 = 5'hd == pms_2 ? io_in_13_Re : _GEN_132; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_134 = 5'he == pms_2 ? io_in_14_Re : _GEN_133; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_135 = 5'hf == pms_2 ? io_in_15_Re : _GEN_134; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_136 = 5'h10 == pms_2 ? io_in_16_Re : _GEN_135; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_137 = 5'h11 == pms_2 ? io_in_17_Re : _GEN_136; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_138 = 5'h12 == pms_2 ? io_in_18_Re : _GEN_137; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_139 = 5'h13 == pms_2 ? io_in_19_Re : _GEN_138; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_140 = 5'h14 == pms_2 ? io_in_20_Re : _GEN_139; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_141 = 5'h15 == pms_2 ? io_in_21_Re : _GEN_140; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_142 = 5'h16 == pms_2 ? io_in_22_Re : _GEN_141; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_145 = 5'h1 == pms_3 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_146 = 5'h2 == pms_3 ? io_in_2_Im : _GEN_145; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_147 = 5'h3 == pms_3 ? io_in_3_Im : _GEN_146; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_148 = 5'h4 == pms_3 ? io_in_4_Im : _GEN_147; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_149 = 5'h5 == pms_3 ? io_in_5_Im : _GEN_148; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_150 = 5'h6 == pms_3 ? io_in_6_Im : _GEN_149; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_151 = 5'h7 == pms_3 ? io_in_7_Im : _GEN_150; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_152 = 5'h8 == pms_3 ? io_in_8_Im : _GEN_151; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_153 = 5'h9 == pms_3 ? io_in_9_Im : _GEN_152; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_154 = 5'ha == pms_3 ? io_in_10_Im : _GEN_153; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_155 = 5'hb == pms_3 ? io_in_11_Im : _GEN_154; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_156 = 5'hc == pms_3 ? io_in_12_Im : _GEN_155; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_157 = 5'hd == pms_3 ? io_in_13_Im : _GEN_156; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_158 = 5'he == pms_3 ? io_in_14_Im : _GEN_157; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_159 = 5'hf == pms_3 ? io_in_15_Im : _GEN_158; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_160 = 5'h10 == pms_3 ? io_in_16_Im : _GEN_159; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_161 = 5'h11 == pms_3 ? io_in_17_Im : _GEN_160; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_162 = 5'h12 == pms_3 ? io_in_18_Im : _GEN_161; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_163 = 5'h13 == pms_3 ? io_in_19_Im : _GEN_162; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_164 = 5'h14 == pms_3 ? io_in_20_Im : _GEN_163; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_165 = 5'h15 == pms_3 ? io_in_21_Im : _GEN_164; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_166 = 5'h16 == pms_3 ? io_in_22_Im : _GEN_165; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_169 = 5'h1 == pms_3 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_170 = 5'h2 == pms_3 ? io_in_2_Re : _GEN_169; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_171 = 5'h3 == pms_3 ? io_in_3_Re : _GEN_170; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_172 = 5'h4 == pms_3 ? io_in_4_Re : _GEN_171; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_173 = 5'h5 == pms_3 ? io_in_5_Re : _GEN_172; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_174 = 5'h6 == pms_3 ? io_in_6_Re : _GEN_173; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_175 = 5'h7 == pms_3 ? io_in_7_Re : _GEN_174; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_176 = 5'h8 == pms_3 ? io_in_8_Re : _GEN_175; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_177 = 5'h9 == pms_3 ? io_in_9_Re : _GEN_176; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_178 = 5'ha == pms_3 ? io_in_10_Re : _GEN_177; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_179 = 5'hb == pms_3 ? io_in_11_Re : _GEN_178; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_180 = 5'hc == pms_3 ? io_in_12_Re : _GEN_179; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_181 = 5'hd == pms_3 ? io_in_13_Re : _GEN_180; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_182 = 5'he == pms_3 ? io_in_14_Re : _GEN_181; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_183 = 5'hf == pms_3 ? io_in_15_Re : _GEN_182; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_184 = 5'h10 == pms_3 ? io_in_16_Re : _GEN_183; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_185 = 5'h11 == pms_3 ? io_in_17_Re : _GEN_184; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_186 = 5'h12 == pms_3 ? io_in_18_Re : _GEN_185; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_187 = 5'h13 == pms_3 ? io_in_19_Re : _GEN_186; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_188 = 5'h14 == pms_3 ? io_in_20_Re : _GEN_187; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_189 = 5'h15 == pms_3 ? io_in_21_Re : _GEN_188; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_190 = 5'h16 == pms_3 ? io_in_22_Re : _GEN_189; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_193 = 5'h1 == pms_4 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_194 = 5'h2 == pms_4 ? io_in_2_Im : _GEN_193; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_195 = 5'h3 == pms_4 ? io_in_3_Im : _GEN_194; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_196 = 5'h4 == pms_4 ? io_in_4_Im : _GEN_195; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_197 = 5'h5 == pms_4 ? io_in_5_Im : _GEN_196; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_198 = 5'h6 == pms_4 ? io_in_6_Im : _GEN_197; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_199 = 5'h7 == pms_4 ? io_in_7_Im : _GEN_198; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_200 = 5'h8 == pms_4 ? io_in_8_Im : _GEN_199; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_201 = 5'h9 == pms_4 ? io_in_9_Im : _GEN_200; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_202 = 5'ha == pms_4 ? io_in_10_Im : _GEN_201; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_203 = 5'hb == pms_4 ? io_in_11_Im : _GEN_202; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_204 = 5'hc == pms_4 ? io_in_12_Im : _GEN_203; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_205 = 5'hd == pms_4 ? io_in_13_Im : _GEN_204; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_206 = 5'he == pms_4 ? io_in_14_Im : _GEN_205; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_207 = 5'hf == pms_4 ? io_in_15_Im : _GEN_206; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_208 = 5'h10 == pms_4 ? io_in_16_Im : _GEN_207; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_209 = 5'h11 == pms_4 ? io_in_17_Im : _GEN_208; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_210 = 5'h12 == pms_4 ? io_in_18_Im : _GEN_209; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_211 = 5'h13 == pms_4 ? io_in_19_Im : _GEN_210; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_212 = 5'h14 == pms_4 ? io_in_20_Im : _GEN_211; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_213 = 5'h15 == pms_4 ? io_in_21_Im : _GEN_212; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_214 = 5'h16 == pms_4 ? io_in_22_Im : _GEN_213; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_217 = 5'h1 == pms_4 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_218 = 5'h2 == pms_4 ? io_in_2_Re : _GEN_217; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_219 = 5'h3 == pms_4 ? io_in_3_Re : _GEN_218; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_220 = 5'h4 == pms_4 ? io_in_4_Re : _GEN_219; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_221 = 5'h5 == pms_4 ? io_in_5_Re : _GEN_220; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_222 = 5'h6 == pms_4 ? io_in_6_Re : _GEN_221; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_223 = 5'h7 == pms_4 ? io_in_7_Re : _GEN_222; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_224 = 5'h8 == pms_4 ? io_in_8_Re : _GEN_223; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_225 = 5'h9 == pms_4 ? io_in_9_Re : _GEN_224; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_226 = 5'ha == pms_4 ? io_in_10_Re : _GEN_225; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_227 = 5'hb == pms_4 ? io_in_11_Re : _GEN_226; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_228 = 5'hc == pms_4 ? io_in_12_Re : _GEN_227; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_229 = 5'hd == pms_4 ? io_in_13_Re : _GEN_228; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_230 = 5'he == pms_4 ? io_in_14_Re : _GEN_229; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_231 = 5'hf == pms_4 ? io_in_15_Re : _GEN_230; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_232 = 5'h10 == pms_4 ? io_in_16_Re : _GEN_231; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_233 = 5'h11 == pms_4 ? io_in_17_Re : _GEN_232; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_234 = 5'h12 == pms_4 ? io_in_18_Re : _GEN_233; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_235 = 5'h13 == pms_4 ? io_in_19_Re : _GEN_234; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_236 = 5'h14 == pms_4 ? io_in_20_Re : _GEN_235; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_237 = 5'h15 == pms_4 ? io_in_21_Re : _GEN_236; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_238 = 5'h16 == pms_4 ? io_in_22_Re : _GEN_237; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_241 = 5'h1 == pms_5 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_242 = 5'h2 == pms_5 ? io_in_2_Im : _GEN_241; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_243 = 5'h3 == pms_5 ? io_in_3_Im : _GEN_242; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_244 = 5'h4 == pms_5 ? io_in_4_Im : _GEN_243; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_245 = 5'h5 == pms_5 ? io_in_5_Im : _GEN_244; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_246 = 5'h6 == pms_5 ? io_in_6_Im : _GEN_245; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_247 = 5'h7 == pms_5 ? io_in_7_Im : _GEN_246; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_248 = 5'h8 == pms_5 ? io_in_8_Im : _GEN_247; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_249 = 5'h9 == pms_5 ? io_in_9_Im : _GEN_248; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_250 = 5'ha == pms_5 ? io_in_10_Im : _GEN_249; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_251 = 5'hb == pms_5 ? io_in_11_Im : _GEN_250; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_252 = 5'hc == pms_5 ? io_in_12_Im : _GEN_251; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_253 = 5'hd == pms_5 ? io_in_13_Im : _GEN_252; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_254 = 5'he == pms_5 ? io_in_14_Im : _GEN_253; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_255 = 5'hf == pms_5 ? io_in_15_Im : _GEN_254; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_256 = 5'h10 == pms_5 ? io_in_16_Im : _GEN_255; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_257 = 5'h11 == pms_5 ? io_in_17_Im : _GEN_256; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_258 = 5'h12 == pms_5 ? io_in_18_Im : _GEN_257; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_259 = 5'h13 == pms_5 ? io_in_19_Im : _GEN_258; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_260 = 5'h14 == pms_5 ? io_in_20_Im : _GEN_259; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_261 = 5'h15 == pms_5 ? io_in_21_Im : _GEN_260; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_262 = 5'h16 == pms_5 ? io_in_22_Im : _GEN_261; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_265 = 5'h1 == pms_5 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_266 = 5'h2 == pms_5 ? io_in_2_Re : _GEN_265; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_267 = 5'h3 == pms_5 ? io_in_3_Re : _GEN_266; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_268 = 5'h4 == pms_5 ? io_in_4_Re : _GEN_267; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_269 = 5'h5 == pms_5 ? io_in_5_Re : _GEN_268; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_270 = 5'h6 == pms_5 ? io_in_6_Re : _GEN_269; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_271 = 5'h7 == pms_5 ? io_in_7_Re : _GEN_270; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_272 = 5'h8 == pms_5 ? io_in_8_Re : _GEN_271; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_273 = 5'h9 == pms_5 ? io_in_9_Re : _GEN_272; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_274 = 5'ha == pms_5 ? io_in_10_Re : _GEN_273; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_275 = 5'hb == pms_5 ? io_in_11_Re : _GEN_274; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_276 = 5'hc == pms_5 ? io_in_12_Re : _GEN_275; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_277 = 5'hd == pms_5 ? io_in_13_Re : _GEN_276; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_278 = 5'he == pms_5 ? io_in_14_Re : _GEN_277; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_279 = 5'hf == pms_5 ? io_in_15_Re : _GEN_278; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_280 = 5'h10 == pms_5 ? io_in_16_Re : _GEN_279; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_281 = 5'h11 == pms_5 ? io_in_17_Re : _GEN_280; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_282 = 5'h12 == pms_5 ? io_in_18_Re : _GEN_281; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_283 = 5'h13 == pms_5 ? io_in_19_Re : _GEN_282; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_284 = 5'h14 == pms_5 ? io_in_20_Re : _GEN_283; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_285 = 5'h15 == pms_5 ? io_in_21_Re : _GEN_284; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_286 = 5'h16 == pms_5 ? io_in_22_Re : _GEN_285; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_289 = 5'h1 == pms_6 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_290 = 5'h2 == pms_6 ? io_in_2_Im : _GEN_289; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_291 = 5'h3 == pms_6 ? io_in_3_Im : _GEN_290; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_292 = 5'h4 == pms_6 ? io_in_4_Im : _GEN_291; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_293 = 5'h5 == pms_6 ? io_in_5_Im : _GEN_292; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_294 = 5'h6 == pms_6 ? io_in_6_Im : _GEN_293; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_295 = 5'h7 == pms_6 ? io_in_7_Im : _GEN_294; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_296 = 5'h8 == pms_6 ? io_in_8_Im : _GEN_295; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_297 = 5'h9 == pms_6 ? io_in_9_Im : _GEN_296; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_298 = 5'ha == pms_6 ? io_in_10_Im : _GEN_297; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_299 = 5'hb == pms_6 ? io_in_11_Im : _GEN_298; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_300 = 5'hc == pms_6 ? io_in_12_Im : _GEN_299; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_301 = 5'hd == pms_6 ? io_in_13_Im : _GEN_300; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_302 = 5'he == pms_6 ? io_in_14_Im : _GEN_301; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_303 = 5'hf == pms_6 ? io_in_15_Im : _GEN_302; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_304 = 5'h10 == pms_6 ? io_in_16_Im : _GEN_303; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_305 = 5'h11 == pms_6 ? io_in_17_Im : _GEN_304; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_306 = 5'h12 == pms_6 ? io_in_18_Im : _GEN_305; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_307 = 5'h13 == pms_6 ? io_in_19_Im : _GEN_306; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_308 = 5'h14 == pms_6 ? io_in_20_Im : _GEN_307; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_309 = 5'h15 == pms_6 ? io_in_21_Im : _GEN_308; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_310 = 5'h16 == pms_6 ? io_in_22_Im : _GEN_309; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_313 = 5'h1 == pms_6 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_314 = 5'h2 == pms_6 ? io_in_2_Re : _GEN_313; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_315 = 5'h3 == pms_6 ? io_in_3_Re : _GEN_314; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_316 = 5'h4 == pms_6 ? io_in_4_Re : _GEN_315; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_317 = 5'h5 == pms_6 ? io_in_5_Re : _GEN_316; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_318 = 5'h6 == pms_6 ? io_in_6_Re : _GEN_317; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_319 = 5'h7 == pms_6 ? io_in_7_Re : _GEN_318; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_320 = 5'h8 == pms_6 ? io_in_8_Re : _GEN_319; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_321 = 5'h9 == pms_6 ? io_in_9_Re : _GEN_320; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_322 = 5'ha == pms_6 ? io_in_10_Re : _GEN_321; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_323 = 5'hb == pms_6 ? io_in_11_Re : _GEN_322; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_324 = 5'hc == pms_6 ? io_in_12_Re : _GEN_323; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_325 = 5'hd == pms_6 ? io_in_13_Re : _GEN_324; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_326 = 5'he == pms_6 ? io_in_14_Re : _GEN_325; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_327 = 5'hf == pms_6 ? io_in_15_Re : _GEN_326; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_328 = 5'h10 == pms_6 ? io_in_16_Re : _GEN_327; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_329 = 5'h11 == pms_6 ? io_in_17_Re : _GEN_328; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_330 = 5'h12 == pms_6 ? io_in_18_Re : _GEN_329; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_331 = 5'h13 == pms_6 ? io_in_19_Re : _GEN_330; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_332 = 5'h14 == pms_6 ? io_in_20_Re : _GEN_331; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_333 = 5'h15 == pms_6 ? io_in_21_Re : _GEN_332; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_334 = 5'h16 == pms_6 ? io_in_22_Re : _GEN_333; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_337 = 5'h1 == pms_7 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_338 = 5'h2 == pms_7 ? io_in_2_Im : _GEN_337; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_339 = 5'h3 == pms_7 ? io_in_3_Im : _GEN_338; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_340 = 5'h4 == pms_7 ? io_in_4_Im : _GEN_339; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_341 = 5'h5 == pms_7 ? io_in_5_Im : _GEN_340; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_342 = 5'h6 == pms_7 ? io_in_6_Im : _GEN_341; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_343 = 5'h7 == pms_7 ? io_in_7_Im : _GEN_342; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_344 = 5'h8 == pms_7 ? io_in_8_Im : _GEN_343; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_345 = 5'h9 == pms_7 ? io_in_9_Im : _GEN_344; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_346 = 5'ha == pms_7 ? io_in_10_Im : _GEN_345; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_347 = 5'hb == pms_7 ? io_in_11_Im : _GEN_346; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_348 = 5'hc == pms_7 ? io_in_12_Im : _GEN_347; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_349 = 5'hd == pms_7 ? io_in_13_Im : _GEN_348; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_350 = 5'he == pms_7 ? io_in_14_Im : _GEN_349; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_351 = 5'hf == pms_7 ? io_in_15_Im : _GEN_350; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_352 = 5'h10 == pms_7 ? io_in_16_Im : _GEN_351; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_353 = 5'h11 == pms_7 ? io_in_17_Im : _GEN_352; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_354 = 5'h12 == pms_7 ? io_in_18_Im : _GEN_353; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_355 = 5'h13 == pms_7 ? io_in_19_Im : _GEN_354; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_356 = 5'h14 == pms_7 ? io_in_20_Im : _GEN_355; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_357 = 5'h15 == pms_7 ? io_in_21_Im : _GEN_356; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_358 = 5'h16 == pms_7 ? io_in_22_Im : _GEN_357; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_361 = 5'h1 == pms_7 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_362 = 5'h2 == pms_7 ? io_in_2_Re : _GEN_361; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_363 = 5'h3 == pms_7 ? io_in_3_Re : _GEN_362; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_364 = 5'h4 == pms_7 ? io_in_4_Re : _GEN_363; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_365 = 5'h5 == pms_7 ? io_in_5_Re : _GEN_364; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_366 = 5'h6 == pms_7 ? io_in_6_Re : _GEN_365; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_367 = 5'h7 == pms_7 ? io_in_7_Re : _GEN_366; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_368 = 5'h8 == pms_7 ? io_in_8_Re : _GEN_367; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_369 = 5'h9 == pms_7 ? io_in_9_Re : _GEN_368; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_370 = 5'ha == pms_7 ? io_in_10_Re : _GEN_369; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_371 = 5'hb == pms_7 ? io_in_11_Re : _GEN_370; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_372 = 5'hc == pms_7 ? io_in_12_Re : _GEN_371; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_373 = 5'hd == pms_7 ? io_in_13_Re : _GEN_372; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_374 = 5'he == pms_7 ? io_in_14_Re : _GEN_373; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_375 = 5'hf == pms_7 ? io_in_15_Re : _GEN_374; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_376 = 5'h10 == pms_7 ? io_in_16_Re : _GEN_375; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_377 = 5'h11 == pms_7 ? io_in_17_Re : _GEN_376; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_378 = 5'h12 == pms_7 ? io_in_18_Re : _GEN_377; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_379 = 5'h13 == pms_7 ? io_in_19_Re : _GEN_378; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_380 = 5'h14 == pms_7 ? io_in_20_Re : _GEN_379; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_381 = 5'h15 == pms_7 ? io_in_21_Re : _GEN_380; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_382 = 5'h16 == pms_7 ? io_in_22_Re : _GEN_381; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_385 = 5'h1 == pms_8 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_386 = 5'h2 == pms_8 ? io_in_2_Im : _GEN_385; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_387 = 5'h3 == pms_8 ? io_in_3_Im : _GEN_386; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_388 = 5'h4 == pms_8 ? io_in_4_Im : _GEN_387; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_389 = 5'h5 == pms_8 ? io_in_5_Im : _GEN_388; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_390 = 5'h6 == pms_8 ? io_in_6_Im : _GEN_389; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_391 = 5'h7 == pms_8 ? io_in_7_Im : _GEN_390; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_392 = 5'h8 == pms_8 ? io_in_8_Im : _GEN_391; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_393 = 5'h9 == pms_8 ? io_in_9_Im : _GEN_392; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_394 = 5'ha == pms_8 ? io_in_10_Im : _GEN_393; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_395 = 5'hb == pms_8 ? io_in_11_Im : _GEN_394; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_396 = 5'hc == pms_8 ? io_in_12_Im : _GEN_395; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_397 = 5'hd == pms_8 ? io_in_13_Im : _GEN_396; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_398 = 5'he == pms_8 ? io_in_14_Im : _GEN_397; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_399 = 5'hf == pms_8 ? io_in_15_Im : _GEN_398; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_400 = 5'h10 == pms_8 ? io_in_16_Im : _GEN_399; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_401 = 5'h11 == pms_8 ? io_in_17_Im : _GEN_400; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_402 = 5'h12 == pms_8 ? io_in_18_Im : _GEN_401; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_403 = 5'h13 == pms_8 ? io_in_19_Im : _GEN_402; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_404 = 5'h14 == pms_8 ? io_in_20_Im : _GEN_403; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_405 = 5'h15 == pms_8 ? io_in_21_Im : _GEN_404; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_406 = 5'h16 == pms_8 ? io_in_22_Im : _GEN_405; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_409 = 5'h1 == pms_8 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_410 = 5'h2 == pms_8 ? io_in_2_Re : _GEN_409; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_411 = 5'h3 == pms_8 ? io_in_3_Re : _GEN_410; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_412 = 5'h4 == pms_8 ? io_in_4_Re : _GEN_411; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_413 = 5'h5 == pms_8 ? io_in_5_Re : _GEN_412; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_414 = 5'h6 == pms_8 ? io_in_6_Re : _GEN_413; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_415 = 5'h7 == pms_8 ? io_in_7_Re : _GEN_414; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_416 = 5'h8 == pms_8 ? io_in_8_Re : _GEN_415; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_417 = 5'h9 == pms_8 ? io_in_9_Re : _GEN_416; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_418 = 5'ha == pms_8 ? io_in_10_Re : _GEN_417; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_419 = 5'hb == pms_8 ? io_in_11_Re : _GEN_418; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_420 = 5'hc == pms_8 ? io_in_12_Re : _GEN_419; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_421 = 5'hd == pms_8 ? io_in_13_Re : _GEN_420; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_422 = 5'he == pms_8 ? io_in_14_Re : _GEN_421; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_423 = 5'hf == pms_8 ? io_in_15_Re : _GEN_422; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_424 = 5'h10 == pms_8 ? io_in_16_Re : _GEN_423; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_425 = 5'h11 == pms_8 ? io_in_17_Re : _GEN_424; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_426 = 5'h12 == pms_8 ? io_in_18_Re : _GEN_425; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_427 = 5'h13 == pms_8 ? io_in_19_Re : _GEN_426; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_428 = 5'h14 == pms_8 ? io_in_20_Re : _GEN_427; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_429 = 5'h15 == pms_8 ? io_in_21_Re : _GEN_428; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_430 = 5'h16 == pms_8 ? io_in_22_Re : _GEN_429; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_433 = 5'h1 == pms_9 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_434 = 5'h2 == pms_9 ? io_in_2_Im : _GEN_433; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_435 = 5'h3 == pms_9 ? io_in_3_Im : _GEN_434; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_436 = 5'h4 == pms_9 ? io_in_4_Im : _GEN_435; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_437 = 5'h5 == pms_9 ? io_in_5_Im : _GEN_436; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_438 = 5'h6 == pms_9 ? io_in_6_Im : _GEN_437; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_439 = 5'h7 == pms_9 ? io_in_7_Im : _GEN_438; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_440 = 5'h8 == pms_9 ? io_in_8_Im : _GEN_439; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_441 = 5'h9 == pms_9 ? io_in_9_Im : _GEN_440; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_442 = 5'ha == pms_9 ? io_in_10_Im : _GEN_441; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_443 = 5'hb == pms_9 ? io_in_11_Im : _GEN_442; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_444 = 5'hc == pms_9 ? io_in_12_Im : _GEN_443; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_445 = 5'hd == pms_9 ? io_in_13_Im : _GEN_444; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_446 = 5'he == pms_9 ? io_in_14_Im : _GEN_445; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_447 = 5'hf == pms_9 ? io_in_15_Im : _GEN_446; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_448 = 5'h10 == pms_9 ? io_in_16_Im : _GEN_447; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_449 = 5'h11 == pms_9 ? io_in_17_Im : _GEN_448; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_450 = 5'h12 == pms_9 ? io_in_18_Im : _GEN_449; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_451 = 5'h13 == pms_9 ? io_in_19_Im : _GEN_450; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_452 = 5'h14 == pms_9 ? io_in_20_Im : _GEN_451; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_453 = 5'h15 == pms_9 ? io_in_21_Im : _GEN_452; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_454 = 5'h16 == pms_9 ? io_in_22_Im : _GEN_453; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_457 = 5'h1 == pms_9 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_458 = 5'h2 == pms_9 ? io_in_2_Re : _GEN_457; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_459 = 5'h3 == pms_9 ? io_in_3_Re : _GEN_458; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_460 = 5'h4 == pms_9 ? io_in_4_Re : _GEN_459; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_461 = 5'h5 == pms_9 ? io_in_5_Re : _GEN_460; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_462 = 5'h6 == pms_9 ? io_in_6_Re : _GEN_461; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_463 = 5'h7 == pms_9 ? io_in_7_Re : _GEN_462; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_464 = 5'h8 == pms_9 ? io_in_8_Re : _GEN_463; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_465 = 5'h9 == pms_9 ? io_in_9_Re : _GEN_464; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_466 = 5'ha == pms_9 ? io_in_10_Re : _GEN_465; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_467 = 5'hb == pms_9 ? io_in_11_Re : _GEN_466; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_468 = 5'hc == pms_9 ? io_in_12_Re : _GEN_467; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_469 = 5'hd == pms_9 ? io_in_13_Re : _GEN_468; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_470 = 5'he == pms_9 ? io_in_14_Re : _GEN_469; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_471 = 5'hf == pms_9 ? io_in_15_Re : _GEN_470; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_472 = 5'h10 == pms_9 ? io_in_16_Re : _GEN_471; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_473 = 5'h11 == pms_9 ? io_in_17_Re : _GEN_472; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_474 = 5'h12 == pms_9 ? io_in_18_Re : _GEN_473; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_475 = 5'h13 == pms_9 ? io_in_19_Re : _GEN_474; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_476 = 5'h14 == pms_9 ? io_in_20_Re : _GEN_475; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_477 = 5'h15 == pms_9 ? io_in_21_Re : _GEN_476; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_478 = 5'h16 == pms_9 ? io_in_22_Re : _GEN_477; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_481 = 5'h1 == pms_10 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_482 = 5'h2 == pms_10 ? io_in_2_Im : _GEN_481; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_483 = 5'h3 == pms_10 ? io_in_3_Im : _GEN_482; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_484 = 5'h4 == pms_10 ? io_in_4_Im : _GEN_483; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_485 = 5'h5 == pms_10 ? io_in_5_Im : _GEN_484; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_486 = 5'h6 == pms_10 ? io_in_6_Im : _GEN_485; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_487 = 5'h7 == pms_10 ? io_in_7_Im : _GEN_486; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_488 = 5'h8 == pms_10 ? io_in_8_Im : _GEN_487; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_489 = 5'h9 == pms_10 ? io_in_9_Im : _GEN_488; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_490 = 5'ha == pms_10 ? io_in_10_Im : _GEN_489; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_491 = 5'hb == pms_10 ? io_in_11_Im : _GEN_490; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_492 = 5'hc == pms_10 ? io_in_12_Im : _GEN_491; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_493 = 5'hd == pms_10 ? io_in_13_Im : _GEN_492; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_494 = 5'he == pms_10 ? io_in_14_Im : _GEN_493; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_495 = 5'hf == pms_10 ? io_in_15_Im : _GEN_494; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_496 = 5'h10 == pms_10 ? io_in_16_Im : _GEN_495; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_497 = 5'h11 == pms_10 ? io_in_17_Im : _GEN_496; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_498 = 5'h12 == pms_10 ? io_in_18_Im : _GEN_497; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_499 = 5'h13 == pms_10 ? io_in_19_Im : _GEN_498; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_500 = 5'h14 == pms_10 ? io_in_20_Im : _GEN_499; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_501 = 5'h15 == pms_10 ? io_in_21_Im : _GEN_500; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_502 = 5'h16 == pms_10 ? io_in_22_Im : _GEN_501; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_505 = 5'h1 == pms_10 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_506 = 5'h2 == pms_10 ? io_in_2_Re : _GEN_505; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_507 = 5'h3 == pms_10 ? io_in_3_Re : _GEN_506; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_508 = 5'h4 == pms_10 ? io_in_4_Re : _GEN_507; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_509 = 5'h5 == pms_10 ? io_in_5_Re : _GEN_508; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_510 = 5'h6 == pms_10 ? io_in_6_Re : _GEN_509; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_511 = 5'h7 == pms_10 ? io_in_7_Re : _GEN_510; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_512 = 5'h8 == pms_10 ? io_in_8_Re : _GEN_511; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_513 = 5'h9 == pms_10 ? io_in_9_Re : _GEN_512; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_514 = 5'ha == pms_10 ? io_in_10_Re : _GEN_513; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_515 = 5'hb == pms_10 ? io_in_11_Re : _GEN_514; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_516 = 5'hc == pms_10 ? io_in_12_Re : _GEN_515; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_517 = 5'hd == pms_10 ? io_in_13_Re : _GEN_516; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_518 = 5'he == pms_10 ? io_in_14_Re : _GEN_517; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_519 = 5'hf == pms_10 ? io_in_15_Re : _GEN_518; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_520 = 5'h10 == pms_10 ? io_in_16_Re : _GEN_519; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_521 = 5'h11 == pms_10 ? io_in_17_Re : _GEN_520; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_522 = 5'h12 == pms_10 ? io_in_18_Re : _GEN_521; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_523 = 5'h13 == pms_10 ? io_in_19_Re : _GEN_522; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_524 = 5'h14 == pms_10 ? io_in_20_Re : _GEN_523; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_525 = 5'h15 == pms_10 ? io_in_21_Re : _GEN_524; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_526 = 5'h16 == pms_10 ? io_in_22_Re : _GEN_525; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_529 = 5'h1 == pms_11 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_530 = 5'h2 == pms_11 ? io_in_2_Im : _GEN_529; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_531 = 5'h3 == pms_11 ? io_in_3_Im : _GEN_530; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_532 = 5'h4 == pms_11 ? io_in_4_Im : _GEN_531; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_533 = 5'h5 == pms_11 ? io_in_5_Im : _GEN_532; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_534 = 5'h6 == pms_11 ? io_in_6_Im : _GEN_533; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_535 = 5'h7 == pms_11 ? io_in_7_Im : _GEN_534; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_536 = 5'h8 == pms_11 ? io_in_8_Im : _GEN_535; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_537 = 5'h9 == pms_11 ? io_in_9_Im : _GEN_536; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_538 = 5'ha == pms_11 ? io_in_10_Im : _GEN_537; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_539 = 5'hb == pms_11 ? io_in_11_Im : _GEN_538; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_540 = 5'hc == pms_11 ? io_in_12_Im : _GEN_539; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_541 = 5'hd == pms_11 ? io_in_13_Im : _GEN_540; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_542 = 5'he == pms_11 ? io_in_14_Im : _GEN_541; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_543 = 5'hf == pms_11 ? io_in_15_Im : _GEN_542; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_544 = 5'h10 == pms_11 ? io_in_16_Im : _GEN_543; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_545 = 5'h11 == pms_11 ? io_in_17_Im : _GEN_544; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_546 = 5'h12 == pms_11 ? io_in_18_Im : _GEN_545; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_547 = 5'h13 == pms_11 ? io_in_19_Im : _GEN_546; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_548 = 5'h14 == pms_11 ? io_in_20_Im : _GEN_547; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_549 = 5'h15 == pms_11 ? io_in_21_Im : _GEN_548; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_550 = 5'h16 == pms_11 ? io_in_22_Im : _GEN_549; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_553 = 5'h1 == pms_11 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_554 = 5'h2 == pms_11 ? io_in_2_Re : _GEN_553; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_555 = 5'h3 == pms_11 ? io_in_3_Re : _GEN_554; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_556 = 5'h4 == pms_11 ? io_in_4_Re : _GEN_555; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_557 = 5'h5 == pms_11 ? io_in_5_Re : _GEN_556; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_558 = 5'h6 == pms_11 ? io_in_6_Re : _GEN_557; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_559 = 5'h7 == pms_11 ? io_in_7_Re : _GEN_558; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_560 = 5'h8 == pms_11 ? io_in_8_Re : _GEN_559; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_561 = 5'h9 == pms_11 ? io_in_9_Re : _GEN_560; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_562 = 5'ha == pms_11 ? io_in_10_Re : _GEN_561; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_563 = 5'hb == pms_11 ? io_in_11_Re : _GEN_562; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_564 = 5'hc == pms_11 ? io_in_12_Re : _GEN_563; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_565 = 5'hd == pms_11 ? io_in_13_Re : _GEN_564; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_566 = 5'he == pms_11 ? io_in_14_Re : _GEN_565; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_567 = 5'hf == pms_11 ? io_in_15_Re : _GEN_566; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_568 = 5'h10 == pms_11 ? io_in_16_Re : _GEN_567; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_569 = 5'h11 == pms_11 ? io_in_17_Re : _GEN_568; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_570 = 5'h12 == pms_11 ? io_in_18_Re : _GEN_569; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_571 = 5'h13 == pms_11 ? io_in_19_Re : _GEN_570; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_572 = 5'h14 == pms_11 ? io_in_20_Re : _GEN_571; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_573 = 5'h15 == pms_11 ? io_in_21_Re : _GEN_572; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_574 = 5'h16 == pms_11 ? io_in_22_Re : _GEN_573; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_577 = 5'h1 == pms_12 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_578 = 5'h2 == pms_12 ? io_in_2_Im : _GEN_577; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_579 = 5'h3 == pms_12 ? io_in_3_Im : _GEN_578; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_580 = 5'h4 == pms_12 ? io_in_4_Im : _GEN_579; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_581 = 5'h5 == pms_12 ? io_in_5_Im : _GEN_580; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_582 = 5'h6 == pms_12 ? io_in_6_Im : _GEN_581; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_583 = 5'h7 == pms_12 ? io_in_7_Im : _GEN_582; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_584 = 5'h8 == pms_12 ? io_in_8_Im : _GEN_583; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_585 = 5'h9 == pms_12 ? io_in_9_Im : _GEN_584; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_586 = 5'ha == pms_12 ? io_in_10_Im : _GEN_585; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_587 = 5'hb == pms_12 ? io_in_11_Im : _GEN_586; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_588 = 5'hc == pms_12 ? io_in_12_Im : _GEN_587; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_589 = 5'hd == pms_12 ? io_in_13_Im : _GEN_588; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_590 = 5'he == pms_12 ? io_in_14_Im : _GEN_589; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_591 = 5'hf == pms_12 ? io_in_15_Im : _GEN_590; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_592 = 5'h10 == pms_12 ? io_in_16_Im : _GEN_591; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_593 = 5'h11 == pms_12 ? io_in_17_Im : _GEN_592; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_594 = 5'h12 == pms_12 ? io_in_18_Im : _GEN_593; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_595 = 5'h13 == pms_12 ? io_in_19_Im : _GEN_594; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_596 = 5'h14 == pms_12 ? io_in_20_Im : _GEN_595; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_597 = 5'h15 == pms_12 ? io_in_21_Im : _GEN_596; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_598 = 5'h16 == pms_12 ? io_in_22_Im : _GEN_597; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_601 = 5'h1 == pms_12 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_602 = 5'h2 == pms_12 ? io_in_2_Re : _GEN_601; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_603 = 5'h3 == pms_12 ? io_in_3_Re : _GEN_602; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_604 = 5'h4 == pms_12 ? io_in_4_Re : _GEN_603; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_605 = 5'h5 == pms_12 ? io_in_5_Re : _GEN_604; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_606 = 5'h6 == pms_12 ? io_in_6_Re : _GEN_605; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_607 = 5'h7 == pms_12 ? io_in_7_Re : _GEN_606; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_608 = 5'h8 == pms_12 ? io_in_8_Re : _GEN_607; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_609 = 5'h9 == pms_12 ? io_in_9_Re : _GEN_608; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_610 = 5'ha == pms_12 ? io_in_10_Re : _GEN_609; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_611 = 5'hb == pms_12 ? io_in_11_Re : _GEN_610; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_612 = 5'hc == pms_12 ? io_in_12_Re : _GEN_611; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_613 = 5'hd == pms_12 ? io_in_13_Re : _GEN_612; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_614 = 5'he == pms_12 ? io_in_14_Re : _GEN_613; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_615 = 5'hf == pms_12 ? io_in_15_Re : _GEN_614; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_616 = 5'h10 == pms_12 ? io_in_16_Re : _GEN_615; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_617 = 5'h11 == pms_12 ? io_in_17_Re : _GEN_616; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_618 = 5'h12 == pms_12 ? io_in_18_Re : _GEN_617; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_619 = 5'h13 == pms_12 ? io_in_19_Re : _GEN_618; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_620 = 5'h14 == pms_12 ? io_in_20_Re : _GEN_619; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_621 = 5'h15 == pms_12 ? io_in_21_Re : _GEN_620; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_622 = 5'h16 == pms_12 ? io_in_22_Re : _GEN_621; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_625 = 5'h1 == pms_13 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_626 = 5'h2 == pms_13 ? io_in_2_Im : _GEN_625; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_627 = 5'h3 == pms_13 ? io_in_3_Im : _GEN_626; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_628 = 5'h4 == pms_13 ? io_in_4_Im : _GEN_627; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_629 = 5'h5 == pms_13 ? io_in_5_Im : _GEN_628; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_630 = 5'h6 == pms_13 ? io_in_6_Im : _GEN_629; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_631 = 5'h7 == pms_13 ? io_in_7_Im : _GEN_630; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_632 = 5'h8 == pms_13 ? io_in_8_Im : _GEN_631; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_633 = 5'h9 == pms_13 ? io_in_9_Im : _GEN_632; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_634 = 5'ha == pms_13 ? io_in_10_Im : _GEN_633; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_635 = 5'hb == pms_13 ? io_in_11_Im : _GEN_634; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_636 = 5'hc == pms_13 ? io_in_12_Im : _GEN_635; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_637 = 5'hd == pms_13 ? io_in_13_Im : _GEN_636; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_638 = 5'he == pms_13 ? io_in_14_Im : _GEN_637; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_639 = 5'hf == pms_13 ? io_in_15_Im : _GEN_638; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_640 = 5'h10 == pms_13 ? io_in_16_Im : _GEN_639; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_641 = 5'h11 == pms_13 ? io_in_17_Im : _GEN_640; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_642 = 5'h12 == pms_13 ? io_in_18_Im : _GEN_641; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_643 = 5'h13 == pms_13 ? io_in_19_Im : _GEN_642; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_644 = 5'h14 == pms_13 ? io_in_20_Im : _GEN_643; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_645 = 5'h15 == pms_13 ? io_in_21_Im : _GEN_644; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_646 = 5'h16 == pms_13 ? io_in_22_Im : _GEN_645; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_649 = 5'h1 == pms_13 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_650 = 5'h2 == pms_13 ? io_in_2_Re : _GEN_649; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_651 = 5'h3 == pms_13 ? io_in_3_Re : _GEN_650; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_652 = 5'h4 == pms_13 ? io_in_4_Re : _GEN_651; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_653 = 5'h5 == pms_13 ? io_in_5_Re : _GEN_652; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_654 = 5'h6 == pms_13 ? io_in_6_Re : _GEN_653; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_655 = 5'h7 == pms_13 ? io_in_7_Re : _GEN_654; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_656 = 5'h8 == pms_13 ? io_in_8_Re : _GEN_655; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_657 = 5'h9 == pms_13 ? io_in_9_Re : _GEN_656; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_658 = 5'ha == pms_13 ? io_in_10_Re : _GEN_657; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_659 = 5'hb == pms_13 ? io_in_11_Re : _GEN_658; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_660 = 5'hc == pms_13 ? io_in_12_Re : _GEN_659; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_661 = 5'hd == pms_13 ? io_in_13_Re : _GEN_660; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_662 = 5'he == pms_13 ? io_in_14_Re : _GEN_661; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_663 = 5'hf == pms_13 ? io_in_15_Re : _GEN_662; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_664 = 5'h10 == pms_13 ? io_in_16_Re : _GEN_663; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_665 = 5'h11 == pms_13 ? io_in_17_Re : _GEN_664; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_666 = 5'h12 == pms_13 ? io_in_18_Re : _GEN_665; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_667 = 5'h13 == pms_13 ? io_in_19_Re : _GEN_666; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_668 = 5'h14 == pms_13 ? io_in_20_Re : _GEN_667; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_669 = 5'h15 == pms_13 ? io_in_21_Re : _GEN_668; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_670 = 5'h16 == pms_13 ? io_in_22_Re : _GEN_669; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_673 = 5'h1 == pms_14 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_674 = 5'h2 == pms_14 ? io_in_2_Im : _GEN_673; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_675 = 5'h3 == pms_14 ? io_in_3_Im : _GEN_674; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_676 = 5'h4 == pms_14 ? io_in_4_Im : _GEN_675; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_677 = 5'h5 == pms_14 ? io_in_5_Im : _GEN_676; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_678 = 5'h6 == pms_14 ? io_in_6_Im : _GEN_677; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_679 = 5'h7 == pms_14 ? io_in_7_Im : _GEN_678; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_680 = 5'h8 == pms_14 ? io_in_8_Im : _GEN_679; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_681 = 5'h9 == pms_14 ? io_in_9_Im : _GEN_680; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_682 = 5'ha == pms_14 ? io_in_10_Im : _GEN_681; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_683 = 5'hb == pms_14 ? io_in_11_Im : _GEN_682; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_684 = 5'hc == pms_14 ? io_in_12_Im : _GEN_683; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_685 = 5'hd == pms_14 ? io_in_13_Im : _GEN_684; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_686 = 5'he == pms_14 ? io_in_14_Im : _GEN_685; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_687 = 5'hf == pms_14 ? io_in_15_Im : _GEN_686; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_688 = 5'h10 == pms_14 ? io_in_16_Im : _GEN_687; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_689 = 5'h11 == pms_14 ? io_in_17_Im : _GEN_688; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_690 = 5'h12 == pms_14 ? io_in_18_Im : _GEN_689; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_691 = 5'h13 == pms_14 ? io_in_19_Im : _GEN_690; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_692 = 5'h14 == pms_14 ? io_in_20_Im : _GEN_691; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_693 = 5'h15 == pms_14 ? io_in_21_Im : _GEN_692; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_694 = 5'h16 == pms_14 ? io_in_22_Im : _GEN_693; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_697 = 5'h1 == pms_14 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_698 = 5'h2 == pms_14 ? io_in_2_Re : _GEN_697; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_699 = 5'h3 == pms_14 ? io_in_3_Re : _GEN_698; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_700 = 5'h4 == pms_14 ? io_in_4_Re : _GEN_699; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_701 = 5'h5 == pms_14 ? io_in_5_Re : _GEN_700; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_702 = 5'h6 == pms_14 ? io_in_6_Re : _GEN_701; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_703 = 5'h7 == pms_14 ? io_in_7_Re : _GEN_702; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_704 = 5'h8 == pms_14 ? io_in_8_Re : _GEN_703; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_705 = 5'h9 == pms_14 ? io_in_9_Re : _GEN_704; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_706 = 5'ha == pms_14 ? io_in_10_Re : _GEN_705; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_707 = 5'hb == pms_14 ? io_in_11_Re : _GEN_706; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_708 = 5'hc == pms_14 ? io_in_12_Re : _GEN_707; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_709 = 5'hd == pms_14 ? io_in_13_Re : _GEN_708; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_710 = 5'he == pms_14 ? io_in_14_Re : _GEN_709; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_711 = 5'hf == pms_14 ? io_in_15_Re : _GEN_710; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_712 = 5'h10 == pms_14 ? io_in_16_Re : _GEN_711; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_713 = 5'h11 == pms_14 ? io_in_17_Re : _GEN_712; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_714 = 5'h12 == pms_14 ? io_in_18_Re : _GEN_713; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_715 = 5'h13 == pms_14 ? io_in_19_Re : _GEN_714; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_716 = 5'h14 == pms_14 ? io_in_20_Re : _GEN_715; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_717 = 5'h15 == pms_14 ? io_in_21_Re : _GEN_716; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_718 = 5'h16 == pms_14 ? io_in_22_Re : _GEN_717; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_721 = 5'h1 == pms_15 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_722 = 5'h2 == pms_15 ? io_in_2_Im : _GEN_721; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_723 = 5'h3 == pms_15 ? io_in_3_Im : _GEN_722; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_724 = 5'h4 == pms_15 ? io_in_4_Im : _GEN_723; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_725 = 5'h5 == pms_15 ? io_in_5_Im : _GEN_724; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_726 = 5'h6 == pms_15 ? io_in_6_Im : _GEN_725; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_727 = 5'h7 == pms_15 ? io_in_7_Im : _GEN_726; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_728 = 5'h8 == pms_15 ? io_in_8_Im : _GEN_727; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_729 = 5'h9 == pms_15 ? io_in_9_Im : _GEN_728; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_730 = 5'ha == pms_15 ? io_in_10_Im : _GEN_729; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_731 = 5'hb == pms_15 ? io_in_11_Im : _GEN_730; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_732 = 5'hc == pms_15 ? io_in_12_Im : _GEN_731; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_733 = 5'hd == pms_15 ? io_in_13_Im : _GEN_732; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_734 = 5'he == pms_15 ? io_in_14_Im : _GEN_733; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_735 = 5'hf == pms_15 ? io_in_15_Im : _GEN_734; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_736 = 5'h10 == pms_15 ? io_in_16_Im : _GEN_735; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_737 = 5'h11 == pms_15 ? io_in_17_Im : _GEN_736; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_738 = 5'h12 == pms_15 ? io_in_18_Im : _GEN_737; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_739 = 5'h13 == pms_15 ? io_in_19_Im : _GEN_738; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_740 = 5'h14 == pms_15 ? io_in_20_Im : _GEN_739; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_741 = 5'h15 == pms_15 ? io_in_21_Im : _GEN_740; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_742 = 5'h16 == pms_15 ? io_in_22_Im : _GEN_741; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_745 = 5'h1 == pms_15 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_746 = 5'h2 == pms_15 ? io_in_2_Re : _GEN_745; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_747 = 5'h3 == pms_15 ? io_in_3_Re : _GEN_746; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_748 = 5'h4 == pms_15 ? io_in_4_Re : _GEN_747; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_749 = 5'h5 == pms_15 ? io_in_5_Re : _GEN_748; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_750 = 5'h6 == pms_15 ? io_in_6_Re : _GEN_749; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_751 = 5'h7 == pms_15 ? io_in_7_Re : _GEN_750; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_752 = 5'h8 == pms_15 ? io_in_8_Re : _GEN_751; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_753 = 5'h9 == pms_15 ? io_in_9_Re : _GEN_752; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_754 = 5'ha == pms_15 ? io_in_10_Re : _GEN_753; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_755 = 5'hb == pms_15 ? io_in_11_Re : _GEN_754; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_756 = 5'hc == pms_15 ? io_in_12_Re : _GEN_755; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_757 = 5'hd == pms_15 ? io_in_13_Re : _GEN_756; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_758 = 5'he == pms_15 ? io_in_14_Re : _GEN_757; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_759 = 5'hf == pms_15 ? io_in_15_Re : _GEN_758; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_760 = 5'h10 == pms_15 ? io_in_16_Re : _GEN_759; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_761 = 5'h11 == pms_15 ? io_in_17_Re : _GEN_760; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_762 = 5'h12 == pms_15 ? io_in_18_Re : _GEN_761; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_763 = 5'h13 == pms_15 ? io_in_19_Re : _GEN_762; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_764 = 5'h14 == pms_15 ? io_in_20_Re : _GEN_763; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_765 = 5'h15 == pms_15 ? io_in_21_Re : _GEN_764; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_766 = 5'h16 == pms_15 ? io_in_22_Re : _GEN_765; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_769 = 5'h1 == pms_16 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_770 = 5'h2 == pms_16 ? io_in_2_Im : _GEN_769; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_771 = 5'h3 == pms_16 ? io_in_3_Im : _GEN_770; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_772 = 5'h4 == pms_16 ? io_in_4_Im : _GEN_771; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_773 = 5'h5 == pms_16 ? io_in_5_Im : _GEN_772; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_774 = 5'h6 == pms_16 ? io_in_6_Im : _GEN_773; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_775 = 5'h7 == pms_16 ? io_in_7_Im : _GEN_774; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_776 = 5'h8 == pms_16 ? io_in_8_Im : _GEN_775; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_777 = 5'h9 == pms_16 ? io_in_9_Im : _GEN_776; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_778 = 5'ha == pms_16 ? io_in_10_Im : _GEN_777; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_779 = 5'hb == pms_16 ? io_in_11_Im : _GEN_778; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_780 = 5'hc == pms_16 ? io_in_12_Im : _GEN_779; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_781 = 5'hd == pms_16 ? io_in_13_Im : _GEN_780; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_782 = 5'he == pms_16 ? io_in_14_Im : _GEN_781; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_783 = 5'hf == pms_16 ? io_in_15_Im : _GEN_782; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_784 = 5'h10 == pms_16 ? io_in_16_Im : _GEN_783; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_785 = 5'h11 == pms_16 ? io_in_17_Im : _GEN_784; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_786 = 5'h12 == pms_16 ? io_in_18_Im : _GEN_785; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_787 = 5'h13 == pms_16 ? io_in_19_Im : _GEN_786; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_788 = 5'h14 == pms_16 ? io_in_20_Im : _GEN_787; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_789 = 5'h15 == pms_16 ? io_in_21_Im : _GEN_788; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_790 = 5'h16 == pms_16 ? io_in_22_Im : _GEN_789; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_793 = 5'h1 == pms_16 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_794 = 5'h2 == pms_16 ? io_in_2_Re : _GEN_793; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_795 = 5'h3 == pms_16 ? io_in_3_Re : _GEN_794; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_796 = 5'h4 == pms_16 ? io_in_4_Re : _GEN_795; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_797 = 5'h5 == pms_16 ? io_in_5_Re : _GEN_796; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_798 = 5'h6 == pms_16 ? io_in_6_Re : _GEN_797; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_799 = 5'h7 == pms_16 ? io_in_7_Re : _GEN_798; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_800 = 5'h8 == pms_16 ? io_in_8_Re : _GEN_799; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_801 = 5'h9 == pms_16 ? io_in_9_Re : _GEN_800; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_802 = 5'ha == pms_16 ? io_in_10_Re : _GEN_801; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_803 = 5'hb == pms_16 ? io_in_11_Re : _GEN_802; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_804 = 5'hc == pms_16 ? io_in_12_Re : _GEN_803; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_805 = 5'hd == pms_16 ? io_in_13_Re : _GEN_804; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_806 = 5'he == pms_16 ? io_in_14_Re : _GEN_805; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_807 = 5'hf == pms_16 ? io_in_15_Re : _GEN_806; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_808 = 5'h10 == pms_16 ? io_in_16_Re : _GEN_807; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_809 = 5'h11 == pms_16 ? io_in_17_Re : _GEN_808; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_810 = 5'h12 == pms_16 ? io_in_18_Re : _GEN_809; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_811 = 5'h13 == pms_16 ? io_in_19_Re : _GEN_810; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_812 = 5'h14 == pms_16 ? io_in_20_Re : _GEN_811; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_813 = 5'h15 == pms_16 ? io_in_21_Re : _GEN_812; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_814 = 5'h16 == pms_16 ? io_in_22_Re : _GEN_813; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_817 = 5'h1 == pms_17 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_818 = 5'h2 == pms_17 ? io_in_2_Im : _GEN_817; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_819 = 5'h3 == pms_17 ? io_in_3_Im : _GEN_818; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_820 = 5'h4 == pms_17 ? io_in_4_Im : _GEN_819; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_821 = 5'h5 == pms_17 ? io_in_5_Im : _GEN_820; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_822 = 5'h6 == pms_17 ? io_in_6_Im : _GEN_821; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_823 = 5'h7 == pms_17 ? io_in_7_Im : _GEN_822; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_824 = 5'h8 == pms_17 ? io_in_8_Im : _GEN_823; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_825 = 5'h9 == pms_17 ? io_in_9_Im : _GEN_824; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_826 = 5'ha == pms_17 ? io_in_10_Im : _GEN_825; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_827 = 5'hb == pms_17 ? io_in_11_Im : _GEN_826; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_828 = 5'hc == pms_17 ? io_in_12_Im : _GEN_827; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_829 = 5'hd == pms_17 ? io_in_13_Im : _GEN_828; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_830 = 5'he == pms_17 ? io_in_14_Im : _GEN_829; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_831 = 5'hf == pms_17 ? io_in_15_Im : _GEN_830; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_832 = 5'h10 == pms_17 ? io_in_16_Im : _GEN_831; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_833 = 5'h11 == pms_17 ? io_in_17_Im : _GEN_832; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_834 = 5'h12 == pms_17 ? io_in_18_Im : _GEN_833; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_835 = 5'h13 == pms_17 ? io_in_19_Im : _GEN_834; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_836 = 5'h14 == pms_17 ? io_in_20_Im : _GEN_835; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_837 = 5'h15 == pms_17 ? io_in_21_Im : _GEN_836; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_838 = 5'h16 == pms_17 ? io_in_22_Im : _GEN_837; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_841 = 5'h1 == pms_17 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_842 = 5'h2 == pms_17 ? io_in_2_Re : _GEN_841; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_843 = 5'h3 == pms_17 ? io_in_3_Re : _GEN_842; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_844 = 5'h4 == pms_17 ? io_in_4_Re : _GEN_843; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_845 = 5'h5 == pms_17 ? io_in_5_Re : _GEN_844; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_846 = 5'h6 == pms_17 ? io_in_6_Re : _GEN_845; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_847 = 5'h7 == pms_17 ? io_in_7_Re : _GEN_846; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_848 = 5'h8 == pms_17 ? io_in_8_Re : _GEN_847; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_849 = 5'h9 == pms_17 ? io_in_9_Re : _GEN_848; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_850 = 5'ha == pms_17 ? io_in_10_Re : _GEN_849; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_851 = 5'hb == pms_17 ? io_in_11_Re : _GEN_850; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_852 = 5'hc == pms_17 ? io_in_12_Re : _GEN_851; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_853 = 5'hd == pms_17 ? io_in_13_Re : _GEN_852; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_854 = 5'he == pms_17 ? io_in_14_Re : _GEN_853; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_855 = 5'hf == pms_17 ? io_in_15_Re : _GEN_854; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_856 = 5'h10 == pms_17 ? io_in_16_Re : _GEN_855; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_857 = 5'h11 == pms_17 ? io_in_17_Re : _GEN_856; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_858 = 5'h12 == pms_17 ? io_in_18_Re : _GEN_857; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_859 = 5'h13 == pms_17 ? io_in_19_Re : _GEN_858; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_860 = 5'h14 == pms_17 ? io_in_20_Re : _GEN_859; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_861 = 5'h15 == pms_17 ? io_in_21_Re : _GEN_860; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_862 = 5'h16 == pms_17 ? io_in_22_Re : _GEN_861; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_865 = 5'h1 == pms_18 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_866 = 5'h2 == pms_18 ? io_in_2_Im : _GEN_865; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_867 = 5'h3 == pms_18 ? io_in_3_Im : _GEN_866; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_868 = 5'h4 == pms_18 ? io_in_4_Im : _GEN_867; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_869 = 5'h5 == pms_18 ? io_in_5_Im : _GEN_868; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_870 = 5'h6 == pms_18 ? io_in_6_Im : _GEN_869; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_871 = 5'h7 == pms_18 ? io_in_7_Im : _GEN_870; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_872 = 5'h8 == pms_18 ? io_in_8_Im : _GEN_871; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_873 = 5'h9 == pms_18 ? io_in_9_Im : _GEN_872; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_874 = 5'ha == pms_18 ? io_in_10_Im : _GEN_873; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_875 = 5'hb == pms_18 ? io_in_11_Im : _GEN_874; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_876 = 5'hc == pms_18 ? io_in_12_Im : _GEN_875; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_877 = 5'hd == pms_18 ? io_in_13_Im : _GEN_876; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_878 = 5'he == pms_18 ? io_in_14_Im : _GEN_877; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_879 = 5'hf == pms_18 ? io_in_15_Im : _GEN_878; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_880 = 5'h10 == pms_18 ? io_in_16_Im : _GEN_879; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_881 = 5'h11 == pms_18 ? io_in_17_Im : _GEN_880; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_882 = 5'h12 == pms_18 ? io_in_18_Im : _GEN_881; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_883 = 5'h13 == pms_18 ? io_in_19_Im : _GEN_882; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_884 = 5'h14 == pms_18 ? io_in_20_Im : _GEN_883; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_885 = 5'h15 == pms_18 ? io_in_21_Im : _GEN_884; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_886 = 5'h16 == pms_18 ? io_in_22_Im : _GEN_885; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_889 = 5'h1 == pms_18 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_890 = 5'h2 == pms_18 ? io_in_2_Re : _GEN_889; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_891 = 5'h3 == pms_18 ? io_in_3_Re : _GEN_890; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_892 = 5'h4 == pms_18 ? io_in_4_Re : _GEN_891; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_893 = 5'h5 == pms_18 ? io_in_5_Re : _GEN_892; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_894 = 5'h6 == pms_18 ? io_in_6_Re : _GEN_893; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_895 = 5'h7 == pms_18 ? io_in_7_Re : _GEN_894; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_896 = 5'h8 == pms_18 ? io_in_8_Re : _GEN_895; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_897 = 5'h9 == pms_18 ? io_in_9_Re : _GEN_896; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_898 = 5'ha == pms_18 ? io_in_10_Re : _GEN_897; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_899 = 5'hb == pms_18 ? io_in_11_Re : _GEN_898; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_900 = 5'hc == pms_18 ? io_in_12_Re : _GEN_899; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_901 = 5'hd == pms_18 ? io_in_13_Re : _GEN_900; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_902 = 5'he == pms_18 ? io_in_14_Re : _GEN_901; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_903 = 5'hf == pms_18 ? io_in_15_Re : _GEN_902; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_904 = 5'h10 == pms_18 ? io_in_16_Re : _GEN_903; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_905 = 5'h11 == pms_18 ? io_in_17_Re : _GEN_904; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_906 = 5'h12 == pms_18 ? io_in_18_Re : _GEN_905; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_907 = 5'h13 == pms_18 ? io_in_19_Re : _GEN_906; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_908 = 5'h14 == pms_18 ? io_in_20_Re : _GEN_907; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_909 = 5'h15 == pms_18 ? io_in_21_Re : _GEN_908; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_910 = 5'h16 == pms_18 ? io_in_22_Re : _GEN_909; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_913 = 5'h1 == pms_19 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_914 = 5'h2 == pms_19 ? io_in_2_Im : _GEN_913; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_915 = 5'h3 == pms_19 ? io_in_3_Im : _GEN_914; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_916 = 5'h4 == pms_19 ? io_in_4_Im : _GEN_915; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_917 = 5'h5 == pms_19 ? io_in_5_Im : _GEN_916; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_918 = 5'h6 == pms_19 ? io_in_6_Im : _GEN_917; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_919 = 5'h7 == pms_19 ? io_in_7_Im : _GEN_918; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_920 = 5'h8 == pms_19 ? io_in_8_Im : _GEN_919; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_921 = 5'h9 == pms_19 ? io_in_9_Im : _GEN_920; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_922 = 5'ha == pms_19 ? io_in_10_Im : _GEN_921; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_923 = 5'hb == pms_19 ? io_in_11_Im : _GEN_922; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_924 = 5'hc == pms_19 ? io_in_12_Im : _GEN_923; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_925 = 5'hd == pms_19 ? io_in_13_Im : _GEN_924; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_926 = 5'he == pms_19 ? io_in_14_Im : _GEN_925; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_927 = 5'hf == pms_19 ? io_in_15_Im : _GEN_926; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_928 = 5'h10 == pms_19 ? io_in_16_Im : _GEN_927; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_929 = 5'h11 == pms_19 ? io_in_17_Im : _GEN_928; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_930 = 5'h12 == pms_19 ? io_in_18_Im : _GEN_929; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_931 = 5'h13 == pms_19 ? io_in_19_Im : _GEN_930; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_932 = 5'h14 == pms_19 ? io_in_20_Im : _GEN_931; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_933 = 5'h15 == pms_19 ? io_in_21_Im : _GEN_932; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_934 = 5'h16 == pms_19 ? io_in_22_Im : _GEN_933; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_937 = 5'h1 == pms_19 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_938 = 5'h2 == pms_19 ? io_in_2_Re : _GEN_937; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_939 = 5'h3 == pms_19 ? io_in_3_Re : _GEN_938; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_940 = 5'h4 == pms_19 ? io_in_4_Re : _GEN_939; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_941 = 5'h5 == pms_19 ? io_in_5_Re : _GEN_940; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_942 = 5'h6 == pms_19 ? io_in_6_Re : _GEN_941; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_943 = 5'h7 == pms_19 ? io_in_7_Re : _GEN_942; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_944 = 5'h8 == pms_19 ? io_in_8_Re : _GEN_943; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_945 = 5'h9 == pms_19 ? io_in_9_Re : _GEN_944; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_946 = 5'ha == pms_19 ? io_in_10_Re : _GEN_945; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_947 = 5'hb == pms_19 ? io_in_11_Re : _GEN_946; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_948 = 5'hc == pms_19 ? io_in_12_Re : _GEN_947; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_949 = 5'hd == pms_19 ? io_in_13_Re : _GEN_948; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_950 = 5'he == pms_19 ? io_in_14_Re : _GEN_949; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_951 = 5'hf == pms_19 ? io_in_15_Re : _GEN_950; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_952 = 5'h10 == pms_19 ? io_in_16_Re : _GEN_951; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_953 = 5'h11 == pms_19 ? io_in_17_Re : _GEN_952; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_954 = 5'h12 == pms_19 ? io_in_18_Re : _GEN_953; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_955 = 5'h13 == pms_19 ? io_in_19_Re : _GEN_954; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_956 = 5'h14 == pms_19 ? io_in_20_Re : _GEN_955; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_957 = 5'h15 == pms_19 ? io_in_21_Re : _GEN_956; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_958 = 5'h16 == pms_19 ? io_in_22_Re : _GEN_957; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_961 = 5'h1 == pms_20 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_962 = 5'h2 == pms_20 ? io_in_2_Im : _GEN_961; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_963 = 5'h3 == pms_20 ? io_in_3_Im : _GEN_962; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_964 = 5'h4 == pms_20 ? io_in_4_Im : _GEN_963; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_965 = 5'h5 == pms_20 ? io_in_5_Im : _GEN_964; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_966 = 5'h6 == pms_20 ? io_in_6_Im : _GEN_965; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_967 = 5'h7 == pms_20 ? io_in_7_Im : _GEN_966; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_968 = 5'h8 == pms_20 ? io_in_8_Im : _GEN_967; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_969 = 5'h9 == pms_20 ? io_in_9_Im : _GEN_968; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_970 = 5'ha == pms_20 ? io_in_10_Im : _GEN_969; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_971 = 5'hb == pms_20 ? io_in_11_Im : _GEN_970; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_972 = 5'hc == pms_20 ? io_in_12_Im : _GEN_971; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_973 = 5'hd == pms_20 ? io_in_13_Im : _GEN_972; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_974 = 5'he == pms_20 ? io_in_14_Im : _GEN_973; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_975 = 5'hf == pms_20 ? io_in_15_Im : _GEN_974; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_976 = 5'h10 == pms_20 ? io_in_16_Im : _GEN_975; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_977 = 5'h11 == pms_20 ? io_in_17_Im : _GEN_976; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_978 = 5'h12 == pms_20 ? io_in_18_Im : _GEN_977; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_979 = 5'h13 == pms_20 ? io_in_19_Im : _GEN_978; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_980 = 5'h14 == pms_20 ? io_in_20_Im : _GEN_979; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_981 = 5'h15 == pms_20 ? io_in_21_Im : _GEN_980; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_982 = 5'h16 == pms_20 ? io_in_22_Im : _GEN_981; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_985 = 5'h1 == pms_20 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_986 = 5'h2 == pms_20 ? io_in_2_Re : _GEN_985; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_987 = 5'h3 == pms_20 ? io_in_3_Re : _GEN_986; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_988 = 5'h4 == pms_20 ? io_in_4_Re : _GEN_987; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_989 = 5'h5 == pms_20 ? io_in_5_Re : _GEN_988; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_990 = 5'h6 == pms_20 ? io_in_6_Re : _GEN_989; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_991 = 5'h7 == pms_20 ? io_in_7_Re : _GEN_990; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_992 = 5'h8 == pms_20 ? io_in_8_Re : _GEN_991; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_993 = 5'h9 == pms_20 ? io_in_9_Re : _GEN_992; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_994 = 5'ha == pms_20 ? io_in_10_Re : _GEN_993; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_995 = 5'hb == pms_20 ? io_in_11_Re : _GEN_994; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_996 = 5'hc == pms_20 ? io_in_12_Re : _GEN_995; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_997 = 5'hd == pms_20 ? io_in_13_Re : _GEN_996; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_998 = 5'he == pms_20 ? io_in_14_Re : _GEN_997; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_999 = 5'hf == pms_20 ? io_in_15_Re : _GEN_998; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1000 = 5'h10 == pms_20 ? io_in_16_Re : _GEN_999; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1001 = 5'h11 == pms_20 ? io_in_17_Re : _GEN_1000; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1002 = 5'h12 == pms_20 ? io_in_18_Re : _GEN_1001; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1003 = 5'h13 == pms_20 ? io_in_19_Re : _GEN_1002; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1004 = 5'h14 == pms_20 ? io_in_20_Re : _GEN_1003; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1005 = 5'h15 == pms_20 ? io_in_21_Re : _GEN_1004; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1006 = 5'h16 == pms_20 ? io_in_22_Re : _GEN_1005; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1009 = 5'h1 == pms_21 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1010 = 5'h2 == pms_21 ? io_in_2_Im : _GEN_1009; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1011 = 5'h3 == pms_21 ? io_in_3_Im : _GEN_1010; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1012 = 5'h4 == pms_21 ? io_in_4_Im : _GEN_1011; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1013 = 5'h5 == pms_21 ? io_in_5_Im : _GEN_1012; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1014 = 5'h6 == pms_21 ? io_in_6_Im : _GEN_1013; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1015 = 5'h7 == pms_21 ? io_in_7_Im : _GEN_1014; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1016 = 5'h8 == pms_21 ? io_in_8_Im : _GEN_1015; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1017 = 5'h9 == pms_21 ? io_in_9_Im : _GEN_1016; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1018 = 5'ha == pms_21 ? io_in_10_Im : _GEN_1017; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1019 = 5'hb == pms_21 ? io_in_11_Im : _GEN_1018; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1020 = 5'hc == pms_21 ? io_in_12_Im : _GEN_1019; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1021 = 5'hd == pms_21 ? io_in_13_Im : _GEN_1020; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1022 = 5'he == pms_21 ? io_in_14_Im : _GEN_1021; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1023 = 5'hf == pms_21 ? io_in_15_Im : _GEN_1022; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1024 = 5'h10 == pms_21 ? io_in_16_Im : _GEN_1023; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1025 = 5'h11 == pms_21 ? io_in_17_Im : _GEN_1024; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1026 = 5'h12 == pms_21 ? io_in_18_Im : _GEN_1025; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1027 = 5'h13 == pms_21 ? io_in_19_Im : _GEN_1026; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1028 = 5'h14 == pms_21 ? io_in_20_Im : _GEN_1027; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1029 = 5'h15 == pms_21 ? io_in_21_Im : _GEN_1028; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1030 = 5'h16 == pms_21 ? io_in_22_Im : _GEN_1029; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1033 = 5'h1 == pms_21 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1034 = 5'h2 == pms_21 ? io_in_2_Re : _GEN_1033; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1035 = 5'h3 == pms_21 ? io_in_3_Re : _GEN_1034; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1036 = 5'h4 == pms_21 ? io_in_4_Re : _GEN_1035; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1037 = 5'h5 == pms_21 ? io_in_5_Re : _GEN_1036; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1038 = 5'h6 == pms_21 ? io_in_6_Re : _GEN_1037; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1039 = 5'h7 == pms_21 ? io_in_7_Re : _GEN_1038; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1040 = 5'h8 == pms_21 ? io_in_8_Re : _GEN_1039; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1041 = 5'h9 == pms_21 ? io_in_9_Re : _GEN_1040; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1042 = 5'ha == pms_21 ? io_in_10_Re : _GEN_1041; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1043 = 5'hb == pms_21 ? io_in_11_Re : _GEN_1042; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1044 = 5'hc == pms_21 ? io_in_12_Re : _GEN_1043; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1045 = 5'hd == pms_21 ? io_in_13_Re : _GEN_1044; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1046 = 5'he == pms_21 ? io_in_14_Re : _GEN_1045; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1047 = 5'hf == pms_21 ? io_in_15_Re : _GEN_1046; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1048 = 5'h10 == pms_21 ? io_in_16_Re : _GEN_1047; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1049 = 5'h11 == pms_21 ? io_in_17_Re : _GEN_1048; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1050 = 5'h12 == pms_21 ? io_in_18_Re : _GEN_1049; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1051 = 5'h13 == pms_21 ? io_in_19_Re : _GEN_1050; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1052 = 5'h14 == pms_21 ? io_in_20_Re : _GEN_1051; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1053 = 5'h15 == pms_21 ? io_in_21_Re : _GEN_1052; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1054 = 5'h16 == pms_21 ? io_in_22_Re : _GEN_1053; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1057 = 5'h1 == pms_22 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1058 = 5'h2 == pms_22 ? io_in_2_Im : _GEN_1057; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1059 = 5'h3 == pms_22 ? io_in_3_Im : _GEN_1058; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1060 = 5'h4 == pms_22 ? io_in_4_Im : _GEN_1059; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1061 = 5'h5 == pms_22 ? io_in_5_Im : _GEN_1060; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1062 = 5'h6 == pms_22 ? io_in_6_Im : _GEN_1061; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1063 = 5'h7 == pms_22 ? io_in_7_Im : _GEN_1062; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1064 = 5'h8 == pms_22 ? io_in_8_Im : _GEN_1063; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1065 = 5'h9 == pms_22 ? io_in_9_Im : _GEN_1064; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1066 = 5'ha == pms_22 ? io_in_10_Im : _GEN_1065; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1067 = 5'hb == pms_22 ? io_in_11_Im : _GEN_1066; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1068 = 5'hc == pms_22 ? io_in_12_Im : _GEN_1067; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1069 = 5'hd == pms_22 ? io_in_13_Im : _GEN_1068; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1070 = 5'he == pms_22 ? io_in_14_Im : _GEN_1069; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1071 = 5'hf == pms_22 ? io_in_15_Im : _GEN_1070; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1072 = 5'h10 == pms_22 ? io_in_16_Im : _GEN_1071; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1073 = 5'h11 == pms_22 ? io_in_17_Im : _GEN_1072; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1074 = 5'h12 == pms_22 ? io_in_18_Im : _GEN_1073; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1075 = 5'h13 == pms_22 ? io_in_19_Im : _GEN_1074; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1076 = 5'h14 == pms_22 ? io_in_20_Im : _GEN_1075; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1077 = 5'h15 == pms_22 ? io_in_21_Im : _GEN_1076; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1078 = 5'h16 == pms_22 ? io_in_22_Im : _GEN_1077; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1081 = 5'h1 == pms_22 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1082 = 5'h2 == pms_22 ? io_in_2_Re : _GEN_1081; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1083 = 5'h3 == pms_22 ? io_in_3_Re : _GEN_1082; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1084 = 5'h4 == pms_22 ? io_in_4_Re : _GEN_1083; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1085 = 5'h5 == pms_22 ? io_in_5_Re : _GEN_1084; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1086 = 5'h6 == pms_22 ? io_in_6_Re : _GEN_1085; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1087 = 5'h7 == pms_22 ? io_in_7_Re : _GEN_1086; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1088 = 5'h8 == pms_22 ? io_in_8_Re : _GEN_1087; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1089 = 5'h9 == pms_22 ? io_in_9_Re : _GEN_1088; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1090 = 5'ha == pms_22 ? io_in_10_Re : _GEN_1089; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1091 = 5'hb == pms_22 ? io_in_11_Re : _GEN_1090; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1092 = 5'hc == pms_22 ? io_in_12_Re : _GEN_1091; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1093 = 5'hd == pms_22 ? io_in_13_Re : _GEN_1092; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1094 = 5'he == pms_22 ? io_in_14_Re : _GEN_1093; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1095 = 5'hf == pms_22 ? io_in_15_Re : _GEN_1094; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1096 = 5'h10 == pms_22 ? io_in_16_Re : _GEN_1095; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1097 = 5'h11 == pms_22 ? io_in_17_Re : _GEN_1096; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1098 = 5'h12 == pms_22 ? io_in_18_Re : _GEN_1097; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1099 = 5'h13 == pms_22 ? io_in_19_Re : _GEN_1098; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1100 = 5'h14 == pms_22 ? io_in_20_Re : _GEN_1099; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1101 = 5'h15 == pms_22 ? io_in_21_Re : _GEN_1100; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1102 = 5'h16 == pms_22 ? io_in_22_Re : _GEN_1101; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1105 = 5'h1 == pms_23 ? io_in_1_Im : io_in_0_Im; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1106 = 5'h2 == pms_23 ? io_in_2_Im : _GEN_1105; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1107 = 5'h3 == pms_23 ? io_in_3_Im : _GEN_1106; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1108 = 5'h4 == pms_23 ? io_in_4_Im : _GEN_1107; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1109 = 5'h5 == pms_23 ? io_in_5_Im : _GEN_1108; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1110 = 5'h6 == pms_23 ? io_in_6_Im : _GEN_1109; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1111 = 5'h7 == pms_23 ? io_in_7_Im : _GEN_1110; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1112 = 5'h8 == pms_23 ? io_in_8_Im : _GEN_1111; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1113 = 5'h9 == pms_23 ? io_in_9_Im : _GEN_1112; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1114 = 5'ha == pms_23 ? io_in_10_Im : _GEN_1113; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1115 = 5'hb == pms_23 ? io_in_11_Im : _GEN_1114; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1116 = 5'hc == pms_23 ? io_in_12_Im : _GEN_1115; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1117 = 5'hd == pms_23 ? io_in_13_Im : _GEN_1116; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1118 = 5'he == pms_23 ? io_in_14_Im : _GEN_1117; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1119 = 5'hf == pms_23 ? io_in_15_Im : _GEN_1118; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1120 = 5'h10 == pms_23 ? io_in_16_Im : _GEN_1119; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1121 = 5'h11 == pms_23 ? io_in_17_Im : _GEN_1120; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1122 = 5'h12 == pms_23 ? io_in_18_Im : _GEN_1121; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1123 = 5'h13 == pms_23 ? io_in_19_Im : _GEN_1122; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1124 = 5'h14 == pms_23 ? io_in_20_Im : _GEN_1123; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1125 = 5'h15 == pms_23 ? io_in_21_Im : _GEN_1124; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1126 = 5'h16 == pms_23 ? io_in_22_Im : _GEN_1125; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1129 = 5'h1 == pms_23 ? io_in_1_Re : io_in_0_Re; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1130 = 5'h2 == pms_23 ? io_in_2_Re : _GEN_1129; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1131 = 5'h3 == pms_23 ? io_in_3_Re : _GEN_1130; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1132 = 5'h4 == pms_23 ? io_in_4_Re : _GEN_1131; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1133 = 5'h5 == pms_23 ? io_in_5_Re : _GEN_1132; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1134 = 5'h6 == pms_23 ? io_in_6_Re : _GEN_1133; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1135 = 5'h7 == pms_23 ? io_in_7_Re : _GEN_1134; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1136 = 5'h8 == pms_23 ? io_in_8_Re : _GEN_1135; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1137 = 5'h9 == pms_23 ? io_in_9_Re : _GEN_1136; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1138 = 5'ha == pms_23 ? io_in_10_Re : _GEN_1137; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1139 = 5'hb == pms_23 ? io_in_11_Re : _GEN_1138; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1140 = 5'hc == pms_23 ? io_in_12_Re : _GEN_1139; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1141 = 5'hd == pms_23 ? io_in_13_Re : _GEN_1140; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1142 = 5'he == pms_23 ? io_in_14_Re : _GEN_1141; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1143 = 5'hf == pms_23 ? io_in_15_Re : _GEN_1142; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1144 = 5'h10 == pms_23 ? io_in_16_Re : _GEN_1143; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1145 = 5'h11 == pms_23 ? io_in_17_Re : _GEN_1144; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1146 = 5'h12 == pms_23 ? io_in_18_Re : _GEN_1145; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1147 = 5'h13 == pms_23 ? io_in_19_Re : _GEN_1146; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1148 = 5'h14 == pms_23 ? io_in_20_Re : _GEN_1147; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1149 = 5'h15 == pms_23 ? io_in_21_Re : _GEN_1148; // @[FFTDesigns.scala 3203:{17,17}]
  wire [31:0] _GEN_1150 = 5'h16 == pms_23 ? io_in_22_Re : _GEN_1149; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_0_Re = 5'h17 == pms_0 ? io_in_23_Re : _GEN_46; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_0_Im = 5'h17 == pms_0 ? io_in_23_Im : _GEN_22; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_1_Re = 5'h17 == pms_1 ? io_in_23_Re : _GEN_94; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_1_Im = 5'h17 == pms_1 ? io_in_23_Im : _GEN_70; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_2_Re = 5'h17 == pms_2 ? io_in_23_Re : _GEN_142; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_2_Im = 5'h17 == pms_2 ? io_in_23_Im : _GEN_118; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_3_Re = 5'h17 == pms_3 ? io_in_23_Re : _GEN_190; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_3_Im = 5'h17 == pms_3 ? io_in_23_Im : _GEN_166; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_4_Re = 5'h17 == pms_4 ? io_in_23_Re : _GEN_238; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_4_Im = 5'h17 == pms_4 ? io_in_23_Im : _GEN_214; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_5_Re = 5'h17 == pms_5 ? io_in_23_Re : _GEN_286; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_5_Im = 5'h17 == pms_5 ? io_in_23_Im : _GEN_262; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_6_Re = 5'h17 == pms_6 ? io_in_23_Re : _GEN_334; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_6_Im = 5'h17 == pms_6 ? io_in_23_Im : _GEN_310; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_7_Re = 5'h17 == pms_7 ? io_in_23_Re : _GEN_382; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_7_Im = 5'h17 == pms_7 ? io_in_23_Im : _GEN_358; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_8_Re = 5'h17 == pms_8 ? io_in_23_Re : _GEN_430; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_8_Im = 5'h17 == pms_8 ? io_in_23_Im : _GEN_406; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_9_Re = 5'h17 == pms_9 ? io_in_23_Re : _GEN_478; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_9_Im = 5'h17 == pms_9 ? io_in_23_Im : _GEN_454; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_10_Re = 5'h17 == pms_10 ? io_in_23_Re : _GEN_526; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_10_Im = 5'h17 == pms_10 ? io_in_23_Im : _GEN_502; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_11_Re = 5'h17 == pms_11 ? io_in_23_Re : _GEN_574; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_11_Im = 5'h17 == pms_11 ? io_in_23_Im : _GEN_550; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_12_Re = 5'h17 == pms_12 ? io_in_23_Re : _GEN_622; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_12_Im = 5'h17 == pms_12 ? io_in_23_Im : _GEN_598; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_13_Re = 5'h17 == pms_13 ? io_in_23_Re : _GEN_670; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_13_Im = 5'h17 == pms_13 ? io_in_23_Im : _GEN_646; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_14_Re = 5'h17 == pms_14 ? io_in_23_Re : _GEN_718; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_14_Im = 5'h17 == pms_14 ? io_in_23_Im : _GEN_694; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_15_Re = 5'h17 == pms_15 ? io_in_23_Re : _GEN_766; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_15_Im = 5'h17 == pms_15 ? io_in_23_Im : _GEN_742; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_16_Re = 5'h17 == pms_16 ? io_in_23_Re : _GEN_814; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_16_Im = 5'h17 == pms_16 ? io_in_23_Im : _GEN_790; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_17_Re = 5'h17 == pms_17 ? io_in_23_Re : _GEN_862; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_17_Im = 5'h17 == pms_17 ? io_in_23_Im : _GEN_838; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_18_Re = 5'h17 == pms_18 ? io_in_23_Re : _GEN_910; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_18_Im = 5'h17 == pms_18 ? io_in_23_Im : _GEN_886; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_19_Re = 5'h17 == pms_19 ? io_in_23_Re : _GEN_958; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_19_Im = 5'h17 == pms_19 ? io_in_23_Im : _GEN_934; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_20_Re = 5'h17 == pms_20 ? io_in_23_Re : _GEN_1006; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_20_Im = 5'h17 == pms_20 ? io_in_23_Im : _GEN_982; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_21_Re = 5'h17 == pms_21 ? io_in_23_Re : _GEN_1054; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_21_Im = 5'h17 == pms_21 ? io_in_23_Im : _GEN_1030; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_22_Re = 5'h17 == pms_22 ? io_in_23_Re : _GEN_1102; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_22_Im = 5'h17 == pms_22 ? io_in_23_Im : _GEN_1078; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_23_Re = 5'h17 == pms_23 ? io_in_23_Re : _GEN_1150; // @[FFTDesigns.scala 3203:{17,17}]
  assign io_out_23_Im = 5'h17 == pms_23 ? io_in_23_Im : _GEN_1126; // @[FFTDesigns.scala 3203:{17,17}]
endmodule
module M0_Config_ROM_7(
  input  [1:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6,
  output [2:0] io_out_7,
  output [2:0] io_out_8,
  output [2:0] io_out_9,
  output [2:0] io_out_10,
  output [2:0] io_out_11,
  output [2:0] io_out_12,
  output [2:0] io_out_13,
  output [2:0] io_out_14,
  output [2:0] io_out_15,
  output [2:0] io_out_16,
  output [2:0] io_out_17,
  output [2:0] io_out_18,
  output [2:0] io_out_19,
  output [2:0] io_out_20,
  output [2:0] io_out_21,
  output [2:0] io_out_22,
  output [2:0] io_out_23
);
  wire [2:0] _GEN_1 = 2'h1 == io_in_cnt ? 3'h1 : 3'h0; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_cnt ? 3'h2 : _GEN_1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_33 = 2'h1 == io_in_cnt ? 3'h2 : 3'h1; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_34 = 2'h2 == io_in_cnt ? 3'h3 : _GEN_33; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_65 = 2'h1 == io_in_cnt ? 3'h3 : 3'h2; // @[FFTDesigns.scala 3227:{17,17}]
  wire [2:0] _GEN_66 = 2'h2 == io_in_cnt ? 3'h0 : _GEN_65; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_7 = 2'h3 == io_in_cnt ? 3'h3 : _GEN_2; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_8 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_9 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_10 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_11 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_12 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_13 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_14 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_15 = 2'h3 == io_in_cnt ? 3'h0 : _GEN_34; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_16 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_17 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_18 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_19 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_20 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_21 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_22 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
  assign io_out_23 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_66; // @[FFTDesigns.scala 3227:{17,17}]
endmodule
module M1_Config_ROM_7(
  input  [1:0] io_in_cnt,
  output [2:0] io_out_0,
  output [2:0] io_out_1,
  output [2:0] io_out_2,
  output [2:0] io_out_3,
  output [2:0] io_out_4,
  output [2:0] io_out_5,
  output [2:0] io_out_6,
  output [2:0] io_out_7,
  output [2:0] io_out_8,
  output [2:0] io_out_9,
  output [2:0] io_out_10,
  output [2:0] io_out_11,
  output [2:0] io_out_12,
  output [2:0] io_out_13,
  output [2:0] io_out_14,
  output [2:0] io_out_15,
  output [2:0] io_out_16,
  output [2:0] io_out_17,
  output [2:0] io_out_18,
  output [2:0] io_out_19,
  output [2:0] io_out_20,
  output [2:0] io_out_21,
  output [2:0] io_out_22,
  output [2:0] io_out_23
);
  wire [2:0] _GEN_1 = 2'h1 == io_in_cnt ? 3'h3 : 3'h0; // @[FFTDesigns.scala 3250:{17,17}]
  wire [2:0] _GEN_2 = 2'h2 == io_in_cnt ? 3'h2 : _GEN_1; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_7 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_8 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_9 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_10 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_11 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_12 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_13 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_14 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_15 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_16 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_17 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_18 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_19 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_20 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_21 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_22 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
  assign io_out_23 = 2'h3 == io_in_cnt ? 3'h1 : _GEN_2; // @[FFTDesigns.scala 3250:{17,17}]
endmodule
module Streaming_Permute_Config_7(
  input  [1:0] io_in_cnt,
  output [4:0] io_out_0,
  output [4:0] io_out_1,
  output [4:0] io_out_2,
  output [4:0] io_out_3,
  output [4:0] io_out_4,
  output [4:0] io_out_5,
  output [4:0] io_out_6,
  output [4:0] io_out_7,
  output [4:0] io_out_8,
  output [4:0] io_out_9,
  output [4:0] io_out_10,
  output [4:0] io_out_11,
  output [4:0] io_out_12,
  output [4:0] io_out_13,
  output [4:0] io_out_14,
  output [4:0] io_out_15,
  output [4:0] io_out_16,
  output [4:0] io_out_17,
  output [4:0] io_out_18,
  output [4:0] io_out_19,
  output [4:0] io_out_20,
  output [4:0] io_out_21,
  output [4:0] io_out_22
);
  wire [4:0] _GEN_2 = 2'h2 == io_in_cnt ? 5'h1 : 5'h0; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_6 = 2'h2 == io_in_cnt ? 5'h4 : 5'h3; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_10 = 2'h2 == io_in_cnt ? 5'h7 : 5'h6; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_14 = 2'h2 == io_in_cnt ? 5'ha : 5'h9; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_18 = 2'h2 == io_in_cnt ? 5'hd : 5'hc; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_22 = 2'h2 == io_in_cnt ? 5'h10 : 5'hf; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_26 = 2'h2 == io_in_cnt ? 5'h13 : 5'h12; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_30 = 2'h2 == io_in_cnt ? 5'h16 : 5'h15; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_34 = 2'h2 == io_in_cnt ? 5'h2 : 5'h1; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_38 = 2'h2 == io_in_cnt ? 5'h5 : 5'h4; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_42 = 2'h2 == io_in_cnt ? 5'h8 : 5'h7; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_46 = 2'h2 == io_in_cnt ? 5'hb : 5'ha; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_50 = 2'h2 == io_in_cnt ? 5'he : 5'hd; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_54 = 2'h2 == io_in_cnt ? 5'h11 : 5'h10; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_58 = 2'h2 == io_in_cnt ? 5'h14 : 5'h13; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_62 = 2'h2 == io_in_cnt ? 5'h17 : 5'h16; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_66 = 2'h2 == io_in_cnt ? 5'h0 : 5'h2; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_70 = 2'h2 == io_in_cnt ? 5'h3 : 5'h5; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_74 = 2'h2 == io_in_cnt ? 5'h6 : 5'h8; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_78 = 2'h2 == io_in_cnt ? 5'h9 : 5'hb; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_82 = 2'h2 == io_in_cnt ? 5'hc : 5'he; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_86 = 2'h2 == io_in_cnt ? 5'hf : 5'h11; // @[FFTDesigns.scala 3273:{17,17}]
  wire [4:0] _GEN_90 = 2'h2 == io_in_cnt ? 5'h12 : 5'h14; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_0 = 2'h3 == io_in_cnt ? 5'h2 : _GEN_2; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_1 = 2'h3 == io_in_cnt ? 5'h5 : _GEN_6; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_2 = 2'h3 == io_in_cnt ? 5'h8 : _GEN_10; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_3 = 2'h3 == io_in_cnt ? 5'hb : _GEN_14; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_4 = 2'h3 == io_in_cnt ? 5'he : _GEN_18; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_5 = 2'h3 == io_in_cnt ? 5'h11 : _GEN_22; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_6 = 2'h3 == io_in_cnt ? 5'h14 : _GEN_26; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_7 = 2'h3 == io_in_cnt ? 5'h17 : _GEN_30; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_8 = 2'h3 == io_in_cnt ? 5'h0 : _GEN_34; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_9 = 2'h3 == io_in_cnt ? 5'h3 : _GEN_38; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_10 = 2'h3 == io_in_cnt ? 5'h6 : _GEN_42; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_11 = 2'h3 == io_in_cnt ? 5'h9 : _GEN_46; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_12 = 2'h3 == io_in_cnt ? 5'hc : _GEN_50; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_13 = 2'h3 == io_in_cnt ? 5'hf : _GEN_54; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_14 = 2'h3 == io_in_cnt ? 5'h12 : _GEN_58; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_15 = 2'h3 == io_in_cnt ? 5'h15 : _GEN_62; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_16 = 2'h3 == io_in_cnt ? 5'h1 : _GEN_66; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_17 = 2'h3 == io_in_cnt ? 5'h4 : _GEN_70; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_18 = 2'h3 == io_in_cnt ? 5'h7 : _GEN_74; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_19 = 2'h3 == io_in_cnt ? 5'ha : _GEN_78; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_20 = 2'h3 == io_in_cnt ? 5'hd : _GEN_82; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_21 = 2'h3 == io_in_cnt ? 5'h10 : _GEN_86; // @[FFTDesigns.scala 3273:{17,17}]
  assign io_out_22 = 2'h3 == io_in_cnt ? 5'h13 : _GEN_90; // @[FFTDesigns.scala 3273:{17,17}]
endmodule
module PermutationsWithStreaming_mr(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  input         io_in_en_5,
  input         io_in_en_6,
  input         io_in_en_7,
  input         io_in_en_8,
  input         io_in_en_9,
  input         io_in_en_10,
  input         io_in_en_11,
  input         io_in_en_12,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_16_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_16_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_16_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_16_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_16_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_16_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_16_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_16_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_17_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_17_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_17_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_17_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_17_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_17_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_17_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_17_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_18_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_18_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_18_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_18_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_18_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_18_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_18_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_18_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_19_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_19_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_19_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_19_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_19_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_19_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_19_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_19_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_20_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_20_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_20_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_20_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_20_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_20_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_20_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_20_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_21_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_21_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_21_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_21_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_21_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_21_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_21_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_21_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_22_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_22_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_22_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_22_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_22_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_22_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_22_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_22_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_23_clock; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_23_io_in_raddr; // @[FFTDesigns.scala 2713:26]
  wire [2:0] RAM_Block_23_io_in_waddr; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_23_io_in_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_23_io_in_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_23_io_re; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_23_io_wr; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_23_io_en; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2713:26]
  wire [31:0] RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2713:26]
  wire  RAM_Block_24_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_24_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_24_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_24_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_24_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_24_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_24_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_24_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_24_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_24_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_25_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_25_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_25_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_25_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_25_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_25_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_25_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_25_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_25_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_25_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_26_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_26_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_26_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_26_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_26_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_26_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_26_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_26_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_26_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_26_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_27_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_27_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_27_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_27_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_27_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_27_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_27_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_27_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_27_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_27_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_28_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_28_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_28_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_28_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_28_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_28_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_28_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_28_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_28_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_28_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_29_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_29_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_29_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_29_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_29_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_29_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_29_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_29_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_29_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_29_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_30_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_30_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_30_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_30_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_30_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_30_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_30_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_30_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_30_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_30_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_31_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_31_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_31_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_31_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_31_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_31_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_31_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_31_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_31_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_31_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_32_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_32_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_32_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_32_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_32_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_32_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_32_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_32_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_32_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_32_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_33_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_33_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_33_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_33_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_33_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_33_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_33_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_33_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_33_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_33_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_34_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_34_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_34_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_34_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_34_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_34_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_34_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_34_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_34_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_34_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_35_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_35_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_35_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_35_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_35_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_35_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_35_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_35_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_35_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_35_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_36_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_36_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_36_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_36_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_36_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_36_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_36_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_36_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_36_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_36_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_37_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_37_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_37_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_37_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_37_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_37_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_37_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_37_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_37_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_37_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_38_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_38_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_38_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_38_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_38_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_38_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_38_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_38_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_38_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_38_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_39_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_39_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_39_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_39_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_39_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_39_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_39_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_39_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_39_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_39_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_40_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_40_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_40_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_40_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_40_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_40_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_40_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_40_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_40_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_40_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_41_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_41_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_41_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_41_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_41_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_41_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_41_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_41_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_41_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_41_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_42_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_42_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_42_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_42_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_42_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_42_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_42_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_42_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_42_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_42_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_43_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_43_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_43_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_43_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_43_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_43_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_43_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_43_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_43_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_43_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_44_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_44_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_44_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_44_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_44_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_44_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_44_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_44_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_44_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_44_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_45_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_45_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_45_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_45_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_45_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_45_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_45_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_45_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_45_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_45_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_46_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_46_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_46_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_46_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_46_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_46_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_46_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_46_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_46_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_46_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_47_clock; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_47_io_in_raddr; // @[FFTDesigns.scala 2717:26]
  wire [2:0] RAM_Block_47_io_in_waddr; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_47_io_in_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_47_io_in_data_Im; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_47_io_re; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_47_io_wr; // @[FFTDesigns.scala 2717:26]
  wire  RAM_Block_47_io_en; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_47_io_out_data_Re; // @[FFTDesigns.scala 2717:26]
  wire [31:0] RAM_Block_47_io_out_data_Im; // @[FFTDesigns.scala 2717:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_8_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_8_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_9_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_9_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_10_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_10_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_11_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_11_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_12_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_12_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_13_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_13_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_14_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_14_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_15_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_15_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_16_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_16_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_17_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_17_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_18_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_18_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_19_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_19_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_20_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_20_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_21_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_21_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_22_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_22_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_23_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_in_23_Im; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_7; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_8; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_9; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_10; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_11; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_12; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_13; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_14; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_15; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_16; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_17; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_18; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_19; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_20; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_21; // @[FFTDesigns.scala 2750:28]
  wire [4:0] PermutationModuleStreamed_io_in_config_22; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_16_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_16_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_17_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_17_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_18_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_18_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_19_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_19_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_20_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_20_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_21_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_21_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_22_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_22_Im; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_23_Re; // @[FFTDesigns.scala 2750:28]
  wire [31:0] PermutationModuleStreamed_io_out_23_Im; // @[FFTDesigns.scala 2750:28]
  wire [1:0] M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_8; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_9; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_10; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_11; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_12; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_13; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_14; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_15; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_16; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_17; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_18; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_19; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_20; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_21; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_22; // @[FFTDesigns.scala 2751:29]
  wire [2:0] M0_Config_ROM_io_out_23; // @[FFTDesigns.scala 2751:29]
  wire [1:0] M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_8; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_9; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_10; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_11; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_12; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_13; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_14; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_15; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_16; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_17; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_18; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_19; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_20; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_21; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_22; // @[FFTDesigns.scala 2752:29]
  wire [2:0] M1_Config_ROM_io_out_23; // @[FFTDesigns.scala 2752:29]
  wire [1:0] Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_15; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_16; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_17; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_18; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_19; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_20; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_21; // @[FFTDesigns.scala 2753:31]
  wire [4:0] Streaming_Permute_Config_io_out_22; // @[FFTDesigns.scala 2753:31]
  reg  offset_switch; // @[FFTDesigns.scala 2710:28]
  reg [1:0] cnt2; // @[FFTDesigns.scala 2755:25]
  reg [2:0] cnt; // @[FFTDesigns.scala 2756:24]
  wire [5:0] lo = {io_in_en_5,io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2757:21]
  wire [12:0] _T = {io_in_en_12,io_in_en_11,io_in_en_10,io_in_en_9,io_in_en_8,io_in_en_7,io_in_en_6,lo}; // @[FFTDesigns.scala 2757:21]
  wire  M0_0_re = |_T; // @[FFTDesigns.scala 2757:28]
  wire  _T_2 = cnt2 == 2'h3; // @[FFTDesigns.scala 2758:19]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2761:28]
  wire [2:0] _cnt_T_1 = cnt + 3'h1; // @[FFTDesigns.scala 2764:22]
  wire [1:0] _cnt2_T_1 = cnt2 + 2'h1; // @[FFTDesigns.scala 2767:24]
  wire  _GEN_5 = cnt2 == 2'h3 & cnt == 3'h5 ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2758:69 2761:25]
  wire [3:0] _M0_0_in_raddr_T_1 = 3'h4 * _offset_switch_T; // @[FFTDesigns.scala 2778:56]
  wire [3:0] _GEN_2482 = {{1'd0}, M0_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_0_in_raddr_T_3 = _GEN_2482 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2483 = {{2'd0}, cnt2}; // @[FFTDesigns.scala 2781:34]
  wire [3:0] _M1_0_in_raddr_T_3 = _GEN_2483 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2781:34]
  wire [3:0] _M1_0_in_waddr_T = 3'h4 * offset_switch; // @[FFTDesigns.scala 2782:56]
  wire [3:0] _GEN_2484 = {{1'd0}, M1_Config_ROM_io_out_0}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_0_in_waddr_T_2 = _GEN_2484 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2485 = {{1'd0}, M0_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_1_in_raddr_T_3 = _GEN_2485 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2487 = {{1'd0}, M1_Config_ROM_io_out_1}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_1_in_waddr_T_2 = _GEN_2487 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2488 = {{1'd0}, M0_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_2_in_raddr_T_3 = _GEN_2488 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2490 = {{1'd0}, M1_Config_ROM_io_out_2}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_2_in_waddr_T_2 = _GEN_2490 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2491 = {{1'd0}, M0_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_3_in_raddr_T_3 = _GEN_2491 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2493 = {{1'd0}, M1_Config_ROM_io_out_3}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_3_in_waddr_T_2 = _GEN_2493 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2494 = {{1'd0}, M0_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_4_in_raddr_T_3 = _GEN_2494 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2496 = {{1'd0}, M1_Config_ROM_io_out_4}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_4_in_waddr_T_2 = _GEN_2496 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2497 = {{1'd0}, M0_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_5_in_raddr_T_3 = _GEN_2497 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2499 = {{1'd0}, M1_Config_ROM_io_out_5}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_5_in_waddr_T_2 = _GEN_2499 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2500 = {{1'd0}, M0_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_6_in_raddr_T_3 = _GEN_2500 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2502 = {{1'd0}, M1_Config_ROM_io_out_6}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_6_in_waddr_T_2 = _GEN_2502 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2503 = {{1'd0}, M0_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_7_in_raddr_T_3 = _GEN_2503 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2505 = {{1'd0}, M1_Config_ROM_io_out_7}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_7_in_waddr_T_2 = _GEN_2505 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2506 = {{1'd0}, M0_Config_ROM_io_out_8}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_8_in_raddr_T_3 = _GEN_2506 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2508 = {{1'd0}, M1_Config_ROM_io_out_8}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_8_in_waddr_T_2 = _GEN_2508 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2509 = {{1'd0}, M0_Config_ROM_io_out_9}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_9_in_raddr_T_3 = _GEN_2509 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2511 = {{1'd0}, M1_Config_ROM_io_out_9}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_9_in_waddr_T_2 = _GEN_2511 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2512 = {{1'd0}, M0_Config_ROM_io_out_10}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_10_in_raddr_T_3 = _GEN_2512 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2514 = {{1'd0}, M1_Config_ROM_io_out_10}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_10_in_waddr_T_2 = _GEN_2514 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2515 = {{1'd0}, M0_Config_ROM_io_out_11}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_11_in_raddr_T_3 = _GEN_2515 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2517 = {{1'd0}, M1_Config_ROM_io_out_11}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_11_in_waddr_T_2 = _GEN_2517 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2518 = {{1'd0}, M0_Config_ROM_io_out_12}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_12_in_raddr_T_3 = _GEN_2518 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2520 = {{1'd0}, M1_Config_ROM_io_out_12}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_12_in_waddr_T_2 = _GEN_2520 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2521 = {{1'd0}, M0_Config_ROM_io_out_13}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_13_in_raddr_T_3 = _GEN_2521 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2523 = {{1'd0}, M1_Config_ROM_io_out_13}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_13_in_waddr_T_2 = _GEN_2523 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2524 = {{1'd0}, M0_Config_ROM_io_out_14}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_14_in_raddr_T_3 = _GEN_2524 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2526 = {{1'd0}, M1_Config_ROM_io_out_14}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_14_in_waddr_T_2 = _GEN_2526 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2527 = {{1'd0}, M0_Config_ROM_io_out_15}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_15_in_raddr_T_3 = _GEN_2527 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2529 = {{1'd0}, M1_Config_ROM_io_out_15}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_15_in_waddr_T_2 = _GEN_2529 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2530 = {{1'd0}, M0_Config_ROM_io_out_16}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_16_in_raddr_T_3 = _GEN_2530 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2532 = {{1'd0}, M1_Config_ROM_io_out_16}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_16_in_waddr_T_2 = _GEN_2532 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2533 = {{1'd0}, M0_Config_ROM_io_out_17}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_17_in_raddr_T_3 = _GEN_2533 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2535 = {{1'd0}, M1_Config_ROM_io_out_17}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_17_in_waddr_T_2 = _GEN_2535 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2536 = {{1'd0}, M0_Config_ROM_io_out_18}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_18_in_raddr_T_3 = _GEN_2536 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2538 = {{1'd0}, M1_Config_ROM_io_out_18}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_18_in_waddr_T_2 = _GEN_2538 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2539 = {{1'd0}, M0_Config_ROM_io_out_19}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_19_in_raddr_T_3 = _GEN_2539 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2541 = {{1'd0}, M1_Config_ROM_io_out_19}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_19_in_waddr_T_2 = _GEN_2541 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2542 = {{1'd0}, M0_Config_ROM_io_out_20}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_20_in_raddr_T_3 = _GEN_2542 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2544 = {{1'd0}, M1_Config_ROM_io_out_20}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_20_in_waddr_T_2 = _GEN_2544 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2545 = {{1'd0}, M0_Config_ROM_io_out_21}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_21_in_raddr_T_3 = _GEN_2545 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2547 = {{1'd0}, M1_Config_ROM_io_out_21}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_21_in_waddr_T_2 = _GEN_2547 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2548 = {{1'd0}, M0_Config_ROM_io_out_22}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_22_in_raddr_T_3 = _GEN_2548 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2550 = {{1'd0}, M1_Config_ROM_io_out_22}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_22_in_waddr_T_2 = _GEN_2550 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _GEN_2551 = {{1'd0}, M0_Config_ROM_io_out_23}; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _M0_23_in_raddr_T_3 = _GEN_2551 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2778:46]
  wire [3:0] _GEN_2553 = {{1'd0}, M1_Config_ROM_io_out_23}; // @[FFTDesigns.scala 2782:46]
  wire [3:0] _M1_23_in_waddr_T_2 = _GEN_2553 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2782:46]
  wire [5:0] _GEN_7 = 3'h1 == cnt ? 6'h10 : 6'h0; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_8 = 3'h2 == cnt ? 6'h8 : _GEN_7; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_9 = 3'h3 == cnt ? 6'h0 : _GEN_8; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_10 = 3'h4 == cnt ? 6'h10 : _GEN_9; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_11 = 3'h5 == cnt ? 6'h8 : _GEN_10; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_14 = 3'h2 == cnt ? 4'h1 : 4'h0; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _GEN_15 = 3'h3 == cnt ? 4'h2 : _GEN_14; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _GEN_16 = 3'h4 == cnt ? 4'h2 : _GEN_15; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _GEN_17 = 3'h5 == cnt ? 4'h3 : _GEN_16; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _M0_0_in_waddr_T_2 = _GEN_17 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2799:50]
  wire [3:0] _GEN_19 = _GEN_11 == 6'h0 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_20 = _GEN_11 == 6'h0 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_21 = _GEN_11 == 6'h0 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [5:0] _GEN_24 = 3'h1 == cnt ? 6'h11 : 6'h1; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_25 = 3'h2 == cnt ? 6'h9 : _GEN_24; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_26 = 3'h3 == cnt ? 6'h1 : _GEN_25; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_27 = 3'h4 == cnt ? 6'h11 : _GEN_26; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_28 = 3'h5 == cnt ? 6'h9 : _GEN_27; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_36 = _GEN_28 == 6'h0 ? _M0_0_in_waddr_T_2 : _GEN_19; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_37 = _GEN_28 == 6'h0 ? io_in_1_Im : _GEN_20; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_38 = _GEN_28 == 6'h0 ? io_in_1_Re : _GEN_21; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_41 = 3'h1 == cnt ? 6'h12 : 6'h2; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_42 = 3'h2 == cnt ? 6'ha : _GEN_41; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_43 = 3'h3 == cnt ? 6'h2 : _GEN_42; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_44 = 3'h4 == cnt ? 6'h12 : _GEN_43; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_45 = 3'h5 == cnt ? 6'ha : _GEN_44; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_53 = _GEN_45 == 6'h0 ? _M0_0_in_waddr_T_2 : _GEN_36; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_54 = _GEN_45 == 6'h0 ? io_in_2_Im : _GEN_37; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_55 = _GEN_45 == 6'h0 ? io_in_2_Re : _GEN_38; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_58 = 3'h1 == cnt ? 6'h13 : 6'h3; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_59 = 3'h2 == cnt ? 6'hb : _GEN_58; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_60 = 3'h3 == cnt ? 6'h3 : _GEN_59; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_61 = 3'h4 == cnt ? 6'h13 : _GEN_60; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_62 = 3'h5 == cnt ? 6'hb : _GEN_61; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_70 = _GEN_62 == 6'h0 ? _M0_0_in_waddr_T_2 : _GEN_53; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_71 = _GEN_62 == 6'h0 ? io_in_3_Im : _GEN_54; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_72 = _GEN_62 == 6'h0 ? io_in_3_Re : _GEN_55; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_75 = 3'h1 == cnt ? 6'h14 : 6'h4; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_76 = 3'h2 == cnt ? 6'hc : _GEN_75; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_77 = 3'h3 == cnt ? 6'h4 : _GEN_76; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_78 = 3'h4 == cnt ? 6'h14 : _GEN_77; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_79 = 3'h5 == cnt ? 6'hc : _GEN_78; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_87 = _GEN_79 == 6'h0 ? _M0_0_in_waddr_T_2 : _GEN_70; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_88 = _GEN_79 == 6'h0 ? io_in_4_Im : _GEN_71; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_89 = _GEN_79 == 6'h0 ? io_in_4_Re : _GEN_72; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_92 = 3'h1 == cnt ? 6'h15 : 6'h5; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_93 = 3'h2 == cnt ? 6'hd : _GEN_92; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_94 = 3'h3 == cnt ? 6'h5 : _GEN_93; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_95 = 3'h4 == cnt ? 6'h15 : _GEN_94; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_96 = 3'h5 == cnt ? 6'hd : _GEN_95; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_104 = _GEN_96 == 6'h0 ? _M0_0_in_waddr_T_2 : _GEN_87; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_105 = _GEN_96 == 6'h0 ? io_in_5_Im : _GEN_88; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_106 = _GEN_96 == 6'h0 ? io_in_5_Re : _GEN_89; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_109 = 3'h1 == cnt ? 6'h16 : 6'h6; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_110 = 3'h2 == cnt ? 6'he : _GEN_109; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_111 = 3'h3 == cnt ? 6'h6 : _GEN_110; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_112 = 3'h4 == cnt ? 6'h16 : _GEN_111; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_113 = 3'h5 == cnt ? 6'he : _GEN_112; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_121 = _GEN_113 == 6'h0 ? _M0_0_in_waddr_T_2 : _GEN_104; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_122 = _GEN_113 == 6'h0 ? io_in_6_Im : _GEN_105; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_123 = _GEN_113 == 6'h0 ? io_in_6_Re : _GEN_106; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_126 = 3'h1 == cnt ? 6'h17 : 6'h7; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_127 = 3'h2 == cnt ? 6'hf : _GEN_126; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_128 = 3'h3 == cnt ? 6'h7 : _GEN_127; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_129 = 3'h4 == cnt ? 6'h17 : _GEN_128; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_130 = 3'h5 == cnt ? 6'hf : _GEN_129; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_138 = _GEN_130 == 6'h0 ? _M0_0_in_waddr_T_2 : _GEN_121; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_139 = _GEN_130 == 6'h0 ? io_in_7_Im : _GEN_122; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_140 = _GEN_130 == 6'h0 ? io_in_7_Re : _GEN_123; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_143 = 3'h1 == cnt ? 6'h0 : 6'h8; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_144 = 3'h2 == cnt ? 6'h10 : _GEN_143; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_145 = 3'h3 == cnt ? 6'h8 : _GEN_144; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_146 = 3'h4 == cnt ? 6'h0 : _GEN_145; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_147 = 3'h5 == cnt ? 6'h10 : _GEN_146; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_149 = 3'h1 == cnt ? 4'h1 : 4'h0; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _GEN_150 = 3'h2 == cnt ? 4'h1 : _GEN_149; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _GEN_151 = 3'h3 == cnt ? 4'h2 : _GEN_150; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _GEN_152 = 3'h4 == cnt ? 4'h3 : _GEN_151; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _GEN_153 = 3'h5 == cnt ? 4'h3 : _GEN_152; // @[FFTDesigns.scala 2799:{50,50}]
  wire [3:0] _M0_0_in_waddr_T_26 = _GEN_153 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2799:50]
  wire [3:0] _GEN_155 = _GEN_147 == 6'h0 ? _M0_0_in_waddr_T_26 : _GEN_138; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_156 = _GEN_147 == 6'h0 ? io_in_8_Im : _GEN_139; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_157 = _GEN_147 == 6'h0 ? io_in_8_Re : _GEN_140; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_160 = 3'h1 == cnt ? 6'h1 : 6'h9; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_161 = 3'h2 == cnt ? 6'h11 : _GEN_160; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_162 = 3'h3 == cnt ? 6'h9 : _GEN_161; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_163 = 3'h4 == cnt ? 6'h1 : _GEN_162; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_164 = 3'h5 == cnt ? 6'h11 : _GEN_163; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_172 = _GEN_164 == 6'h0 ? _M0_0_in_waddr_T_26 : _GEN_155; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_173 = _GEN_164 == 6'h0 ? io_in_9_Im : _GEN_156; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_174 = _GEN_164 == 6'h0 ? io_in_9_Re : _GEN_157; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_177 = 3'h1 == cnt ? 6'h2 : 6'ha; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_178 = 3'h2 == cnt ? 6'h12 : _GEN_177; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_179 = 3'h3 == cnt ? 6'ha : _GEN_178; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_180 = 3'h4 == cnt ? 6'h2 : _GEN_179; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_181 = 3'h5 == cnt ? 6'h12 : _GEN_180; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_189 = _GEN_181 == 6'h0 ? _M0_0_in_waddr_T_26 : _GEN_172; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_190 = _GEN_181 == 6'h0 ? io_in_10_Im : _GEN_173; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_191 = _GEN_181 == 6'h0 ? io_in_10_Re : _GEN_174; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_194 = 3'h1 == cnt ? 6'h3 : 6'hb; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_195 = 3'h2 == cnt ? 6'h13 : _GEN_194; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_196 = 3'h3 == cnt ? 6'hb : _GEN_195; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_197 = 3'h4 == cnt ? 6'h3 : _GEN_196; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_198 = 3'h5 == cnt ? 6'h13 : _GEN_197; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_206 = _GEN_198 == 6'h0 ? _M0_0_in_waddr_T_26 : _GEN_189; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_207 = _GEN_198 == 6'h0 ? io_in_11_Im : _GEN_190; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_208 = _GEN_198 == 6'h0 ? io_in_11_Re : _GEN_191; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_211 = 3'h1 == cnt ? 6'h4 : 6'hc; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_212 = 3'h2 == cnt ? 6'h14 : _GEN_211; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_213 = 3'h3 == cnt ? 6'hc : _GEN_212; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_214 = 3'h4 == cnt ? 6'h4 : _GEN_213; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_215 = 3'h5 == cnt ? 6'h14 : _GEN_214; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_223 = _GEN_215 == 6'h0 ? _M0_0_in_waddr_T_26 : _GEN_206; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_224 = _GEN_215 == 6'h0 ? io_in_12_Im : _GEN_207; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_225 = _GEN_215 == 6'h0 ? io_in_12_Re : _GEN_208; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_228 = 3'h1 == cnt ? 6'h5 : 6'hd; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_229 = 3'h2 == cnt ? 6'h15 : _GEN_228; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_230 = 3'h3 == cnt ? 6'hd : _GEN_229; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_231 = 3'h4 == cnt ? 6'h5 : _GEN_230; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_232 = 3'h5 == cnt ? 6'h15 : _GEN_231; // @[FFTDesigns.scala 2797:{35,35}]
  wire [3:0] _GEN_240 = _GEN_232 == 6'h0 ? _M0_0_in_waddr_T_26 : _GEN_223; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_241 = _GEN_232 == 6'h0 ? io_in_13_Im : _GEN_224; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_242 = _GEN_232 == 6'h0 ? io_in_13_Re : _GEN_225; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_245 = 3'h1 == cnt ? 6'h6 : 6'he; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_246 = 3'h2 == cnt ? 6'h16 : _GEN_245; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_247 = 3'h3 == cnt ? 6'he : _GEN_246; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_248 = 3'h4 == cnt ? 6'h6 : _GEN_247; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_249 = 3'h5 == cnt ? 6'h16 : _GEN_248; // @[FFTDesigns.scala 2797:{35,35}]
  wire  _GEN_256 = _GEN_249 == 6'h0 | (_GEN_232 == 6'h0 | (_GEN_215 == 6'h0 | (_GEN_198 == 6'h0 | (_GEN_181 == 6'h0 | (
    _GEN_164 == 6'h0 | (_GEN_147 == 6'h0 | (_GEN_130 == 6'h0 | (_GEN_113 == 6'h0 | (_GEN_96 == 6'h0 | (_GEN_79 == 6'h0
     | (_GEN_62 == 6'h0 | (_GEN_45 == 6'h0 | (_GEN_28 == 6'h0 | _GEN_11 == 6'h0))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_257 = _GEN_249 == 6'h0 ? _M0_0_in_waddr_T_26 : _GEN_240; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_258 = _GEN_249 == 6'h0 ? io_in_14_Im : _GEN_241; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_259 = _GEN_249 == 6'h0 ? io_in_14_Re : _GEN_242; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [5:0] _GEN_262 = 3'h1 == cnt ? 6'h7 : 6'hf; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_263 = 3'h2 == cnt ? 6'h17 : _GEN_262; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_264 = 3'h3 == cnt ? 6'hf : _GEN_263; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_265 = 3'h4 == cnt ? 6'h7 : _GEN_264; // @[FFTDesigns.scala 2797:{35,35}]
  wire [5:0] _GEN_266 = 3'h5 == cnt ? 6'h17 : _GEN_265; // @[FFTDesigns.scala 2797:{35,35}]
  wire  _GEN_273 = _GEN_266 == 6'h0 | _GEN_256; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_274 = _GEN_266 == 6'h0 ? _M0_0_in_waddr_T_26 : _GEN_257; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_275 = _GEN_266 == 6'h0 ? io_in_15_Im : _GEN_258; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_276 = _GEN_266 == 6'h0 ? io_in_15_Re : _GEN_259; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_279 = _GEN_11 == 6'h1 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_280 = _GEN_11 == 6'h1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_281 = _GEN_11 == 6'h1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_284 = _GEN_28 == 6'h1 ? _M0_0_in_waddr_T_2 : _GEN_279; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_285 = _GEN_28 == 6'h1 ? io_in_1_Im : _GEN_280; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_286 = _GEN_28 == 6'h1 ? io_in_1_Re : _GEN_281; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_289 = _GEN_45 == 6'h1 ? _M0_0_in_waddr_T_2 : _GEN_284; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_290 = _GEN_45 == 6'h1 ? io_in_2_Im : _GEN_285; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_291 = _GEN_45 == 6'h1 ? io_in_2_Re : _GEN_286; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_294 = _GEN_62 == 6'h1 ? _M0_0_in_waddr_T_2 : _GEN_289; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_295 = _GEN_62 == 6'h1 ? io_in_3_Im : _GEN_290; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_296 = _GEN_62 == 6'h1 ? io_in_3_Re : _GEN_291; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_299 = _GEN_79 == 6'h1 ? _M0_0_in_waddr_T_2 : _GEN_294; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_300 = _GEN_79 == 6'h1 ? io_in_4_Im : _GEN_295; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_301 = _GEN_79 == 6'h1 ? io_in_4_Re : _GEN_296; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_304 = _GEN_96 == 6'h1 ? _M0_0_in_waddr_T_2 : _GEN_299; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_305 = _GEN_96 == 6'h1 ? io_in_5_Im : _GEN_300; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_306 = _GEN_96 == 6'h1 ? io_in_5_Re : _GEN_301; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_309 = _GEN_113 == 6'h1 ? _M0_0_in_waddr_T_2 : _GEN_304; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_310 = _GEN_113 == 6'h1 ? io_in_6_Im : _GEN_305; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_311 = _GEN_113 == 6'h1 ? io_in_6_Re : _GEN_306; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_314 = _GEN_130 == 6'h1 ? _M0_0_in_waddr_T_2 : _GEN_309; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_315 = _GEN_130 == 6'h1 ? io_in_7_Im : _GEN_310; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_316 = _GEN_130 == 6'h1 ? io_in_7_Re : _GEN_311; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_319 = _GEN_147 == 6'h1 ? _M0_0_in_waddr_T_26 : _GEN_314; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_320 = _GEN_147 == 6'h1 ? io_in_8_Im : _GEN_315; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_321 = _GEN_147 == 6'h1 ? io_in_8_Re : _GEN_316; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_324 = _GEN_164 == 6'h1 ? _M0_0_in_waddr_T_26 : _GEN_319; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_325 = _GEN_164 == 6'h1 ? io_in_9_Im : _GEN_320; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_326 = _GEN_164 == 6'h1 ? io_in_9_Re : _GEN_321; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_329 = _GEN_181 == 6'h1 ? _M0_0_in_waddr_T_26 : _GEN_324; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_330 = _GEN_181 == 6'h1 ? io_in_10_Im : _GEN_325; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_331 = _GEN_181 == 6'h1 ? io_in_10_Re : _GEN_326; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_334 = _GEN_198 == 6'h1 ? _M0_0_in_waddr_T_26 : _GEN_329; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_335 = _GEN_198 == 6'h1 ? io_in_11_Im : _GEN_330; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_336 = _GEN_198 == 6'h1 ? io_in_11_Re : _GEN_331; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_339 = _GEN_215 == 6'h1 ? _M0_0_in_waddr_T_26 : _GEN_334; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_340 = _GEN_215 == 6'h1 ? io_in_12_Im : _GEN_335; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_341 = _GEN_215 == 6'h1 ? io_in_12_Re : _GEN_336; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_344 = _GEN_232 == 6'h1 ? _M0_0_in_waddr_T_26 : _GEN_339; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_345 = _GEN_232 == 6'h1 ? io_in_13_Im : _GEN_340; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_346 = _GEN_232 == 6'h1 ? io_in_13_Re : _GEN_341; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_348 = _GEN_249 == 6'h1 | (_GEN_232 == 6'h1 | (_GEN_215 == 6'h1 | (_GEN_198 == 6'h1 | (_GEN_181 == 6'h1 | (
    _GEN_164 == 6'h1 | (_GEN_147 == 6'h1 | (_GEN_130 == 6'h1 | (_GEN_113 == 6'h1 | (_GEN_96 == 6'h1 | (_GEN_79 == 6'h1
     | (_GEN_62 == 6'h1 | (_GEN_45 == 6'h1 | (_GEN_28 == 6'h1 | _GEN_11 == 6'h1))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_349 = _GEN_249 == 6'h1 ? _M0_0_in_waddr_T_26 : _GEN_344; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_350 = _GEN_249 == 6'h1 ? io_in_14_Im : _GEN_345; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_351 = _GEN_249 == 6'h1 ? io_in_14_Re : _GEN_346; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_353 = _GEN_266 == 6'h1 | _GEN_348; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_354 = _GEN_266 == 6'h1 ? _M0_0_in_waddr_T_26 : _GEN_349; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_355 = _GEN_266 == 6'h1 ? io_in_15_Im : _GEN_350; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_356 = _GEN_266 == 6'h1 ? io_in_15_Re : _GEN_351; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_359 = _GEN_11 == 6'h2 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_360 = _GEN_11 == 6'h2 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_361 = _GEN_11 == 6'h2 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_364 = _GEN_28 == 6'h2 ? _M0_0_in_waddr_T_2 : _GEN_359; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_365 = _GEN_28 == 6'h2 ? io_in_1_Im : _GEN_360; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_366 = _GEN_28 == 6'h2 ? io_in_1_Re : _GEN_361; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_369 = _GEN_45 == 6'h2 ? _M0_0_in_waddr_T_2 : _GEN_364; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_370 = _GEN_45 == 6'h2 ? io_in_2_Im : _GEN_365; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_371 = _GEN_45 == 6'h2 ? io_in_2_Re : _GEN_366; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_374 = _GEN_62 == 6'h2 ? _M0_0_in_waddr_T_2 : _GEN_369; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_375 = _GEN_62 == 6'h2 ? io_in_3_Im : _GEN_370; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_376 = _GEN_62 == 6'h2 ? io_in_3_Re : _GEN_371; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_379 = _GEN_79 == 6'h2 ? _M0_0_in_waddr_T_2 : _GEN_374; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_380 = _GEN_79 == 6'h2 ? io_in_4_Im : _GEN_375; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_381 = _GEN_79 == 6'h2 ? io_in_4_Re : _GEN_376; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_384 = _GEN_96 == 6'h2 ? _M0_0_in_waddr_T_2 : _GEN_379; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_385 = _GEN_96 == 6'h2 ? io_in_5_Im : _GEN_380; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_386 = _GEN_96 == 6'h2 ? io_in_5_Re : _GEN_381; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_389 = _GEN_113 == 6'h2 ? _M0_0_in_waddr_T_2 : _GEN_384; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_390 = _GEN_113 == 6'h2 ? io_in_6_Im : _GEN_385; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_391 = _GEN_113 == 6'h2 ? io_in_6_Re : _GEN_386; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_394 = _GEN_130 == 6'h2 ? _M0_0_in_waddr_T_2 : _GEN_389; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_395 = _GEN_130 == 6'h2 ? io_in_7_Im : _GEN_390; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_396 = _GEN_130 == 6'h2 ? io_in_7_Re : _GEN_391; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_399 = _GEN_147 == 6'h2 ? _M0_0_in_waddr_T_26 : _GEN_394; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_400 = _GEN_147 == 6'h2 ? io_in_8_Im : _GEN_395; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_401 = _GEN_147 == 6'h2 ? io_in_8_Re : _GEN_396; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_404 = _GEN_164 == 6'h2 ? _M0_0_in_waddr_T_26 : _GEN_399; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_405 = _GEN_164 == 6'h2 ? io_in_9_Im : _GEN_400; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_406 = _GEN_164 == 6'h2 ? io_in_9_Re : _GEN_401; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_409 = _GEN_181 == 6'h2 ? _M0_0_in_waddr_T_26 : _GEN_404; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_410 = _GEN_181 == 6'h2 ? io_in_10_Im : _GEN_405; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_411 = _GEN_181 == 6'h2 ? io_in_10_Re : _GEN_406; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_414 = _GEN_198 == 6'h2 ? _M0_0_in_waddr_T_26 : _GEN_409; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_415 = _GEN_198 == 6'h2 ? io_in_11_Im : _GEN_410; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_416 = _GEN_198 == 6'h2 ? io_in_11_Re : _GEN_411; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_419 = _GEN_215 == 6'h2 ? _M0_0_in_waddr_T_26 : _GEN_414; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_420 = _GEN_215 == 6'h2 ? io_in_12_Im : _GEN_415; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_421 = _GEN_215 == 6'h2 ? io_in_12_Re : _GEN_416; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_424 = _GEN_232 == 6'h2 ? _M0_0_in_waddr_T_26 : _GEN_419; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_425 = _GEN_232 == 6'h2 ? io_in_13_Im : _GEN_420; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_426 = _GEN_232 == 6'h2 ? io_in_13_Re : _GEN_421; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_428 = _GEN_249 == 6'h2 | (_GEN_232 == 6'h2 | (_GEN_215 == 6'h2 | (_GEN_198 == 6'h2 | (_GEN_181 == 6'h2 | (
    _GEN_164 == 6'h2 | (_GEN_147 == 6'h2 | (_GEN_130 == 6'h2 | (_GEN_113 == 6'h2 | (_GEN_96 == 6'h2 | (_GEN_79 == 6'h2
     | (_GEN_62 == 6'h2 | (_GEN_45 == 6'h2 | (_GEN_28 == 6'h2 | _GEN_11 == 6'h2))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_429 = _GEN_249 == 6'h2 ? _M0_0_in_waddr_T_26 : _GEN_424; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_430 = _GEN_249 == 6'h2 ? io_in_14_Im : _GEN_425; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_431 = _GEN_249 == 6'h2 ? io_in_14_Re : _GEN_426; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_433 = _GEN_266 == 6'h2 | _GEN_428; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_434 = _GEN_266 == 6'h2 ? _M0_0_in_waddr_T_26 : _GEN_429; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_435 = _GEN_266 == 6'h2 ? io_in_15_Im : _GEN_430; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_436 = _GEN_266 == 6'h2 ? io_in_15_Re : _GEN_431; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_439 = _GEN_11 == 6'h3 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_440 = _GEN_11 == 6'h3 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_441 = _GEN_11 == 6'h3 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_444 = _GEN_28 == 6'h3 ? _M0_0_in_waddr_T_2 : _GEN_439; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_445 = _GEN_28 == 6'h3 ? io_in_1_Im : _GEN_440; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_446 = _GEN_28 == 6'h3 ? io_in_1_Re : _GEN_441; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_449 = _GEN_45 == 6'h3 ? _M0_0_in_waddr_T_2 : _GEN_444; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_450 = _GEN_45 == 6'h3 ? io_in_2_Im : _GEN_445; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_451 = _GEN_45 == 6'h3 ? io_in_2_Re : _GEN_446; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_454 = _GEN_62 == 6'h3 ? _M0_0_in_waddr_T_2 : _GEN_449; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_455 = _GEN_62 == 6'h3 ? io_in_3_Im : _GEN_450; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_456 = _GEN_62 == 6'h3 ? io_in_3_Re : _GEN_451; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_459 = _GEN_79 == 6'h3 ? _M0_0_in_waddr_T_2 : _GEN_454; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_460 = _GEN_79 == 6'h3 ? io_in_4_Im : _GEN_455; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_461 = _GEN_79 == 6'h3 ? io_in_4_Re : _GEN_456; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_464 = _GEN_96 == 6'h3 ? _M0_0_in_waddr_T_2 : _GEN_459; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_465 = _GEN_96 == 6'h3 ? io_in_5_Im : _GEN_460; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_466 = _GEN_96 == 6'h3 ? io_in_5_Re : _GEN_461; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_469 = _GEN_113 == 6'h3 ? _M0_0_in_waddr_T_2 : _GEN_464; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_470 = _GEN_113 == 6'h3 ? io_in_6_Im : _GEN_465; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_471 = _GEN_113 == 6'h3 ? io_in_6_Re : _GEN_466; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_474 = _GEN_130 == 6'h3 ? _M0_0_in_waddr_T_2 : _GEN_469; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_475 = _GEN_130 == 6'h3 ? io_in_7_Im : _GEN_470; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_476 = _GEN_130 == 6'h3 ? io_in_7_Re : _GEN_471; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_479 = _GEN_147 == 6'h3 ? _M0_0_in_waddr_T_26 : _GEN_474; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_480 = _GEN_147 == 6'h3 ? io_in_8_Im : _GEN_475; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_481 = _GEN_147 == 6'h3 ? io_in_8_Re : _GEN_476; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_484 = _GEN_164 == 6'h3 ? _M0_0_in_waddr_T_26 : _GEN_479; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_485 = _GEN_164 == 6'h3 ? io_in_9_Im : _GEN_480; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_486 = _GEN_164 == 6'h3 ? io_in_9_Re : _GEN_481; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_489 = _GEN_181 == 6'h3 ? _M0_0_in_waddr_T_26 : _GEN_484; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_490 = _GEN_181 == 6'h3 ? io_in_10_Im : _GEN_485; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_491 = _GEN_181 == 6'h3 ? io_in_10_Re : _GEN_486; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_494 = _GEN_198 == 6'h3 ? _M0_0_in_waddr_T_26 : _GEN_489; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_495 = _GEN_198 == 6'h3 ? io_in_11_Im : _GEN_490; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_496 = _GEN_198 == 6'h3 ? io_in_11_Re : _GEN_491; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_499 = _GEN_215 == 6'h3 ? _M0_0_in_waddr_T_26 : _GEN_494; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_500 = _GEN_215 == 6'h3 ? io_in_12_Im : _GEN_495; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_501 = _GEN_215 == 6'h3 ? io_in_12_Re : _GEN_496; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_504 = _GEN_232 == 6'h3 ? _M0_0_in_waddr_T_26 : _GEN_499; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_505 = _GEN_232 == 6'h3 ? io_in_13_Im : _GEN_500; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_506 = _GEN_232 == 6'h3 ? io_in_13_Re : _GEN_501; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_508 = _GEN_249 == 6'h3 | (_GEN_232 == 6'h3 | (_GEN_215 == 6'h3 | (_GEN_198 == 6'h3 | (_GEN_181 == 6'h3 | (
    _GEN_164 == 6'h3 | (_GEN_147 == 6'h3 | (_GEN_130 == 6'h3 | (_GEN_113 == 6'h3 | (_GEN_96 == 6'h3 | (_GEN_79 == 6'h3
     | (_GEN_62 == 6'h3 | (_GEN_45 == 6'h3 | (_GEN_28 == 6'h3 | _GEN_11 == 6'h3))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_509 = _GEN_249 == 6'h3 ? _M0_0_in_waddr_T_26 : _GEN_504; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_510 = _GEN_249 == 6'h3 ? io_in_14_Im : _GEN_505; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_511 = _GEN_249 == 6'h3 ? io_in_14_Re : _GEN_506; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_513 = _GEN_266 == 6'h3 | _GEN_508; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_514 = _GEN_266 == 6'h3 ? _M0_0_in_waddr_T_26 : _GEN_509; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_515 = _GEN_266 == 6'h3 ? io_in_15_Im : _GEN_510; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_516 = _GEN_266 == 6'h3 ? io_in_15_Re : _GEN_511; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_519 = _GEN_11 == 6'h4 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_520 = _GEN_11 == 6'h4 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_521 = _GEN_11 == 6'h4 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_524 = _GEN_28 == 6'h4 ? _M0_0_in_waddr_T_2 : _GEN_519; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_525 = _GEN_28 == 6'h4 ? io_in_1_Im : _GEN_520; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_526 = _GEN_28 == 6'h4 ? io_in_1_Re : _GEN_521; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_529 = _GEN_45 == 6'h4 ? _M0_0_in_waddr_T_2 : _GEN_524; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_530 = _GEN_45 == 6'h4 ? io_in_2_Im : _GEN_525; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_531 = _GEN_45 == 6'h4 ? io_in_2_Re : _GEN_526; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_534 = _GEN_62 == 6'h4 ? _M0_0_in_waddr_T_2 : _GEN_529; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_535 = _GEN_62 == 6'h4 ? io_in_3_Im : _GEN_530; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_536 = _GEN_62 == 6'h4 ? io_in_3_Re : _GEN_531; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_539 = _GEN_79 == 6'h4 ? _M0_0_in_waddr_T_2 : _GEN_534; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_540 = _GEN_79 == 6'h4 ? io_in_4_Im : _GEN_535; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_541 = _GEN_79 == 6'h4 ? io_in_4_Re : _GEN_536; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_544 = _GEN_96 == 6'h4 ? _M0_0_in_waddr_T_2 : _GEN_539; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_545 = _GEN_96 == 6'h4 ? io_in_5_Im : _GEN_540; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_546 = _GEN_96 == 6'h4 ? io_in_5_Re : _GEN_541; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_549 = _GEN_113 == 6'h4 ? _M0_0_in_waddr_T_2 : _GEN_544; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_550 = _GEN_113 == 6'h4 ? io_in_6_Im : _GEN_545; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_551 = _GEN_113 == 6'h4 ? io_in_6_Re : _GEN_546; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_554 = _GEN_130 == 6'h4 ? _M0_0_in_waddr_T_2 : _GEN_549; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_555 = _GEN_130 == 6'h4 ? io_in_7_Im : _GEN_550; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_556 = _GEN_130 == 6'h4 ? io_in_7_Re : _GEN_551; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_559 = _GEN_147 == 6'h4 ? _M0_0_in_waddr_T_26 : _GEN_554; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_560 = _GEN_147 == 6'h4 ? io_in_8_Im : _GEN_555; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_561 = _GEN_147 == 6'h4 ? io_in_8_Re : _GEN_556; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_564 = _GEN_164 == 6'h4 ? _M0_0_in_waddr_T_26 : _GEN_559; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_565 = _GEN_164 == 6'h4 ? io_in_9_Im : _GEN_560; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_566 = _GEN_164 == 6'h4 ? io_in_9_Re : _GEN_561; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_569 = _GEN_181 == 6'h4 ? _M0_0_in_waddr_T_26 : _GEN_564; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_570 = _GEN_181 == 6'h4 ? io_in_10_Im : _GEN_565; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_571 = _GEN_181 == 6'h4 ? io_in_10_Re : _GEN_566; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_574 = _GEN_198 == 6'h4 ? _M0_0_in_waddr_T_26 : _GEN_569; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_575 = _GEN_198 == 6'h4 ? io_in_11_Im : _GEN_570; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_576 = _GEN_198 == 6'h4 ? io_in_11_Re : _GEN_571; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_579 = _GEN_215 == 6'h4 ? _M0_0_in_waddr_T_26 : _GEN_574; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_580 = _GEN_215 == 6'h4 ? io_in_12_Im : _GEN_575; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_581 = _GEN_215 == 6'h4 ? io_in_12_Re : _GEN_576; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_584 = _GEN_232 == 6'h4 ? _M0_0_in_waddr_T_26 : _GEN_579; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_585 = _GEN_232 == 6'h4 ? io_in_13_Im : _GEN_580; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_586 = _GEN_232 == 6'h4 ? io_in_13_Re : _GEN_581; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_588 = _GEN_249 == 6'h4 | (_GEN_232 == 6'h4 | (_GEN_215 == 6'h4 | (_GEN_198 == 6'h4 | (_GEN_181 == 6'h4 | (
    _GEN_164 == 6'h4 | (_GEN_147 == 6'h4 | (_GEN_130 == 6'h4 | (_GEN_113 == 6'h4 | (_GEN_96 == 6'h4 | (_GEN_79 == 6'h4
     | (_GEN_62 == 6'h4 | (_GEN_45 == 6'h4 | (_GEN_28 == 6'h4 | _GEN_11 == 6'h4))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_589 = _GEN_249 == 6'h4 ? _M0_0_in_waddr_T_26 : _GEN_584; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_590 = _GEN_249 == 6'h4 ? io_in_14_Im : _GEN_585; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_591 = _GEN_249 == 6'h4 ? io_in_14_Re : _GEN_586; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_593 = _GEN_266 == 6'h4 | _GEN_588; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_594 = _GEN_266 == 6'h4 ? _M0_0_in_waddr_T_26 : _GEN_589; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_595 = _GEN_266 == 6'h4 ? io_in_15_Im : _GEN_590; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_596 = _GEN_266 == 6'h4 ? io_in_15_Re : _GEN_591; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_599 = _GEN_11 == 6'h5 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_600 = _GEN_11 == 6'h5 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_601 = _GEN_11 == 6'h5 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_604 = _GEN_28 == 6'h5 ? _M0_0_in_waddr_T_2 : _GEN_599; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_605 = _GEN_28 == 6'h5 ? io_in_1_Im : _GEN_600; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_606 = _GEN_28 == 6'h5 ? io_in_1_Re : _GEN_601; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_609 = _GEN_45 == 6'h5 ? _M0_0_in_waddr_T_2 : _GEN_604; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_610 = _GEN_45 == 6'h5 ? io_in_2_Im : _GEN_605; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_611 = _GEN_45 == 6'h5 ? io_in_2_Re : _GEN_606; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_614 = _GEN_62 == 6'h5 ? _M0_0_in_waddr_T_2 : _GEN_609; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_615 = _GEN_62 == 6'h5 ? io_in_3_Im : _GEN_610; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_616 = _GEN_62 == 6'h5 ? io_in_3_Re : _GEN_611; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_619 = _GEN_79 == 6'h5 ? _M0_0_in_waddr_T_2 : _GEN_614; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_620 = _GEN_79 == 6'h5 ? io_in_4_Im : _GEN_615; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_621 = _GEN_79 == 6'h5 ? io_in_4_Re : _GEN_616; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_624 = _GEN_96 == 6'h5 ? _M0_0_in_waddr_T_2 : _GEN_619; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_625 = _GEN_96 == 6'h5 ? io_in_5_Im : _GEN_620; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_626 = _GEN_96 == 6'h5 ? io_in_5_Re : _GEN_621; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_629 = _GEN_113 == 6'h5 ? _M0_0_in_waddr_T_2 : _GEN_624; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_630 = _GEN_113 == 6'h5 ? io_in_6_Im : _GEN_625; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_631 = _GEN_113 == 6'h5 ? io_in_6_Re : _GEN_626; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_634 = _GEN_130 == 6'h5 ? _M0_0_in_waddr_T_2 : _GEN_629; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_635 = _GEN_130 == 6'h5 ? io_in_7_Im : _GEN_630; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_636 = _GEN_130 == 6'h5 ? io_in_7_Re : _GEN_631; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_639 = _GEN_147 == 6'h5 ? _M0_0_in_waddr_T_26 : _GEN_634; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_640 = _GEN_147 == 6'h5 ? io_in_8_Im : _GEN_635; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_641 = _GEN_147 == 6'h5 ? io_in_8_Re : _GEN_636; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_644 = _GEN_164 == 6'h5 ? _M0_0_in_waddr_T_26 : _GEN_639; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_645 = _GEN_164 == 6'h5 ? io_in_9_Im : _GEN_640; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_646 = _GEN_164 == 6'h5 ? io_in_9_Re : _GEN_641; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_649 = _GEN_181 == 6'h5 ? _M0_0_in_waddr_T_26 : _GEN_644; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_650 = _GEN_181 == 6'h5 ? io_in_10_Im : _GEN_645; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_651 = _GEN_181 == 6'h5 ? io_in_10_Re : _GEN_646; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_654 = _GEN_198 == 6'h5 ? _M0_0_in_waddr_T_26 : _GEN_649; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_655 = _GEN_198 == 6'h5 ? io_in_11_Im : _GEN_650; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_656 = _GEN_198 == 6'h5 ? io_in_11_Re : _GEN_651; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_659 = _GEN_215 == 6'h5 ? _M0_0_in_waddr_T_26 : _GEN_654; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_660 = _GEN_215 == 6'h5 ? io_in_12_Im : _GEN_655; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_661 = _GEN_215 == 6'h5 ? io_in_12_Re : _GEN_656; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_664 = _GEN_232 == 6'h5 ? _M0_0_in_waddr_T_26 : _GEN_659; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_665 = _GEN_232 == 6'h5 ? io_in_13_Im : _GEN_660; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_666 = _GEN_232 == 6'h5 ? io_in_13_Re : _GEN_661; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_668 = _GEN_249 == 6'h5 | (_GEN_232 == 6'h5 | (_GEN_215 == 6'h5 | (_GEN_198 == 6'h5 | (_GEN_181 == 6'h5 | (
    _GEN_164 == 6'h5 | (_GEN_147 == 6'h5 | (_GEN_130 == 6'h5 | (_GEN_113 == 6'h5 | (_GEN_96 == 6'h5 | (_GEN_79 == 6'h5
     | (_GEN_62 == 6'h5 | (_GEN_45 == 6'h5 | (_GEN_28 == 6'h5 | _GEN_11 == 6'h5))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_669 = _GEN_249 == 6'h5 ? _M0_0_in_waddr_T_26 : _GEN_664; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_670 = _GEN_249 == 6'h5 ? io_in_14_Im : _GEN_665; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_671 = _GEN_249 == 6'h5 ? io_in_14_Re : _GEN_666; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_673 = _GEN_266 == 6'h5 | _GEN_668; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_674 = _GEN_266 == 6'h5 ? _M0_0_in_waddr_T_26 : _GEN_669; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_675 = _GEN_266 == 6'h5 ? io_in_15_Im : _GEN_670; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_676 = _GEN_266 == 6'h5 ? io_in_15_Re : _GEN_671; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_679 = _GEN_11 == 6'h6 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_680 = _GEN_11 == 6'h6 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_681 = _GEN_11 == 6'h6 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_684 = _GEN_28 == 6'h6 ? _M0_0_in_waddr_T_2 : _GEN_679; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_685 = _GEN_28 == 6'h6 ? io_in_1_Im : _GEN_680; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_686 = _GEN_28 == 6'h6 ? io_in_1_Re : _GEN_681; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_689 = _GEN_45 == 6'h6 ? _M0_0_in_waddr_T_2 : _GEN_684; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_690 = _GEN_45 == 6'h6 ? io_in_2_Im : _GEN_685; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_691 = _GEN_45 == 6'h6 ? io_in_2_Re : _GEN_686; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_694 = _GEN_62 == 6'h6 ? _M0_0_in_waddr_T_2 : _GEN_689; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_695 = _GEN_62 == 6'h6 ? io_in_3_Im : _GEN_690; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_696 = _GEN_62 == 6'h6 ? io_in_3_Re : _GEN_691; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_699 = _GEN_79 == 6'h6 ? _M0_0_in_waddr_T_2 : _GEN_694; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_700 = _GEN_79 == 6'h6 ? io_in_4_Im : _GEN_695; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_701 = _GEN_79 == 6'h6 ? io_in_4_Re : _GEN_696; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_704 = _GEN_96 == 6'h6 ? _M0_0_in_waddr_T_2 : _GEN_699; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_705 = _GEN_96 == 6'h6 ? io_in_5_Im : _GEN_700; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_706 = _GEN_96 == 6'h6 ? io_in_5_Re : _GEN_701; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_709 = _GEN_113 == 6'h6 ? _M0_0_in_waddr_T_2 : _GEN_704; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_710 = _GEN_113 == 6'h6 ? io_in_6_Im : _GEN_705; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_711 = _GEN_113 == 6'h6 ? io_in_6_Re : _GEN_706; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_714 = _GEN_130 == 6'h6 ? _M0_0_in_waddr_T_2 : _GEN_709; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_715 = _GEN_130 == 6'h6 ? io_in_7_Im : _GEN_710; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_716 = _GEN_130 == 6'h6 ? io_in_7_Re : _GEN_711; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_719 = _GEN_147 == 6'h6 ? _M0_0_in_waddr_T_26 : _GEN_714; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_720 = _GEN_147 == 6'h6 ? io_in_8_Im : _GEN_715; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_721 = _GEN_147 == 6'h6 ? io_in_8_Re : _GEN_716; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_724 = _GEN_164 == 6'h6 ? _M0_0_in_waddr_T_26 : _GEN_719; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_725 = _GEN_164 == 6'h6 ? io_in_9_Im : _GEN_720; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_726 = _GEN_164 == 6'h6 ? io_in_9_Re : _GEN_721; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_729 = _GEN_181 == 6'h6 ? _M0_0_in_waddr_T_26 : _GEN_724; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_730 = _GEN_181 == 6'h6 ? io_in_10_Im : _GEN_725; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_731 = _GEN_181 == 6'h6 ? io_in_10_Re : _GEN_726; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_734 = _GEN_198 == 6'h6 ? _M0_0_in_waddr_T_26 : _GEN_729; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_735 = _GEN_198 == 6'h6 ? io_in_11_Im : _GEN_730; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_736 = _GEN_198 == 6'h6 ? io_in_11_Re : _GEN_731; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_739 = _GEN_215 == 6'h6 ? _M0_0_in_waddr_T_26 : _GEN_734; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_740 = _GEN_215 == 6'h6 ? io_in_12_Im : _GEN_735; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_741 = _GEN_215 == 6'h6 ? io_in_12_Re : _GEN_736; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_744 = _GEN_232 == 6'h6 ? _M0_0_in_waddr_T_26 : _GEN_739; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_745 = _GEN_232 == 6'h6 ? io_in_13_Im : _GEN_740; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_746 = _GEN_232 == 6'h6 ? io_in_13_Re : _GEN_741; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_748 = _GEN_249 == 6'h6 | (_GEN_232 == 6'h6 | (_GEN_215 == 6'h6 | (_GEN_198 == 6'h6 | (_GEN_181 == 6'h6 | (
    _GEN_164 == 6'h6 | (_GEN_147 == 6'h6 | (_GEN_130 == 6'h6 | (_GEN_113 == 6'h6 | (_GEN_96 == 6'h6 | (_GEN_79 == 6'h6
     | (_GEN_62 == 6'h6 | (_GEN_45 == 6'h6 | (_GEN_28 == 6'h6 | _GEN_11 == 6'h6))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_749 = _GEN_249 == 6'h6 ? _M0_0_in_waddr_T_26 : _GEN_744; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_750 = _GEN_249 == 6'h6 ? io_in_14_Im : _GEN_745; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_751 = _GEN_249 == 6'h6 ? io_in_14_Re : _GEN_746; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_753 = _GEN_266 == 6'h6 | _GEN_748; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_754 = _GEN_266 == 6'h6 ? _M0_0_in_waddr_T_26 : _GEN_749; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_755 = _GEN_266 == 6'h6 ? io_in_15_Im : _GEN_750; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_756 = _GEN_266 == 6'h6 ? io_in_15_Re : _GEN_751; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_759 = _GEN_11 == 6'h7 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_760 = _GEN_11 == 6'h7 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_761 = _GEN_11 == 6'h7 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_764 = _GEN_28 == 6'h7 ? _M0_0_in_waddr_T_2 : _GEN_759; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_765 = _GEN_28 == 6'h7 ? io_in_1_Im : _GEN_760; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_766 = _GEN_28 == 6'h7 ? io_in_1_Re : _GEN_761; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_769 = _GEN_45 == 6'h7 ? _M0_0_in_waddr_T_2 : _GEN_764; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_770 = _GEN_45 == 6'h7 ? io_in_2_Im : _GEN_765; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_771 = _GEN_45 == 6'h7 ? io_in_2_Re : _GEN_766; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_774 = _GEN_62 == 6'h7 ? _M0_0_in_waddr_T_2 : _GEN_769; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_775 = _GEN_62 == 6'h7 ? io_in_3_Im : _GEN_770; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_776 = _GEN_62 == 6'h7 ? io_in_3_Re : _GEN_771; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_779 = _GEN_79 == 6'h7 ? _M0_0_in_waddr_T_2 : _GEN_774; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_780 = _GEN_79 == 6'h7 ? io_in_4_Im : _GEN_775; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_781 = _GEN_79 == 6'h7 ? io_in_4_Re : _GEN_776; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_784 = _GEN_96 == 6'h7 ? _M0_0_in_waddr_T_2 : _GEN_779; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_785 = _GEN_96 == 6'h7 ? io_in_5_Im : _GEN_780; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_786 = _GEN_96 == 6'h7 ? io_in_5_Re : _GEN_781; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_789 = _GEN_113 == 6'h7 ? _M0_0_in_waddr_T_2 : _GEN_784; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_790 = _GEN_113 == 6'h7 ? io_in_6_Im : _GEN_785; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_791 = _GEN_113 == 6'h7 ? io_in_6_Re : _GEN_786; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_794 = _GEN_130 == 6'h7 ? _M0_0_in_waddr_T_2 : _GEN_789; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_795 = _GEN_130 == 6'h7 ? io_in_7_Im : _GEN_790; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_796 = _GEN_130 == 6'h7 ? io_in_7_Re : _GEN_791; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_799 = _GEN_147 == 6'h7 ? _M0_0_in_waddr_T_26 : _GEN_794; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_800 = _GEN_147 == 6'h7 ? io_in_8_Im : _GEN_795; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_801 = _GEN_147 == 6'h7 ? io_in_8_Re : _GEN_796; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_804 = _GEN_164 == 6'h7 ? _M0_0_in_waddr_T_26 : _GEN_799; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_805 = _GEN_164 == 6'h7 ? io_in_9_Im : _GEN_800; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_806 = _GEN_164 == 6'h7 ? io_in_9_Re : _GEN_801; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_809 = _GEN_181 == 6'h7 ? _M0_0_in_waddr_T_26 : _GEN_804; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_810 = _GEN_181 == 6'h7 ? io_in_10_Im : _GEN_805; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_811 = _GEN_181 == 6'h7 ? io_in_10_Re : _GEN_806; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_814 = _GEN_198 == 6'h7 ? _M0_0_in_waddr_T_26 : _GEN_809; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_815 = _GEN_198 == 6'h7 ? io_in_11_Im : _GEN_810; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_816 = _GEN_198 == 6'h7 ? io_in_11_Re : _GEN_811; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_819 = _GEN_215 == 6'h7 ? _M0_0_in_waddr_T_26 : _GEN_814; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_820 = _GEN_215 == 6'h7 ? io_in_12_Im : _GEN_815; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_821 = _GEN_215 == 6'h7 ? io_in_12_Re : _GEN_816; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_824 = _GEN_232 == 6'h7 ? _M0_0_in_waddr_T_26 : _GEN_819; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_825 = _GEN_232 == 6'h7 ? io_in_13_Im : _GEN_820; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_826 = _GEN_232 == 6'h7 ? io_in_13_Re : _GEN_821; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_828 = _GEN_249 == 6'h7 | (_GEN_232 == 6'h7 | (_GEN_215 == 6'h7 | (_GEN_198 == 6'h7 | (_GEN_181 == 6'h7 | (
    _GEN_164 == 6'h7 | (_GEN_147 == 6'h7 | (_GEN_130 == 6'h7 | (_GEN_113 == 6'h7 | (_GEN_96 == 6'h7 | (_GEN_79 == 6'h7
     | (_GEN_62 == 6'h7 | (_GEN_45 == 6'h7 | (_GEN_28 == 6'h7 | _GEN_11 == 6'h7))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_829 = _GEN_249 == 6'h7 ? _M0_0_in_waddr_T_26 : _GEN_824; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_830 = _GEN_249 == 6'h7 ? io_in_14_Im : _GEN_825; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_831 = _GEN_249 == 6'h7 ? io_in_14_Re : _GEN_826; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_833 = _GEN_266 == 6'h7 | _GEN_828; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_834 = _GEN_266 == 6'h7 ? _M0_0_in_waddr_T_26 : _GEN_829; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_835 = _GEN_266 == 6'h7 ? io_in_15_Im : _GEN_830; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_836 = _GEN_266 == 6'h7 ? io_in_15_Re : _GEN_831; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_839 = _GEN_11 == 6'h8 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_840 = _GEN_11 == 6'h8 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_841 = _GEN_11 == 6'h8 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_844 = _GEN_28 == 6'h8 ? _M0_0_in_waddr_T_2 : _GEN_839; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_845 = _GEN_28 == 6'h8 ? io_in_1_Im : _GEN_840; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_846 = _GEN_28 == 6'h8 ? io_in_1_Re : _GEN_841; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_849 = _GEN_45 == 6'h8 ? _M0_0_in_waddr_T_2 : _GEN_844; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_850 = _GEN_45 == 6'h8 ? io_in_2_Im : _GEN_845; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_851 = _GEN_45 == 6'h8 ? io_in_2_Re : _GEN_846; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_854 = _GEN_62 == 6'h8 ? _M0_0_in_waddr_T_2 : _GEN_849; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_855 = _GEN_62 == 6'h8 ? io_in_3_Im : _GEN_850; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_856 = _GEN_62 == 6'h8 ? io_in_3_Re : _GEN_851; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_859 = _GEN_79 == 6'h8 ? _M0_0_in_waddr_T_2 : _GEN_854; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_860 = _GEN_79 == 6'h8 ? io_in_4_Im : _GEN_855; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_861 = _GEN_79 == 6'h8 ? io_in_4_Re : _GEN_856; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_864 = _GEN_96 == 6'h8 ? _M0_0_in_waddr_T_2 : _GEN_859; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_865 = _GEN_96 == 6'h8 ? io_in_5_Im : _GEN_860; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_866 = _GEN_96 == 6'h8 ? io_in_5_Re : _GEN_861; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_869 = _GEN_113 == 6'h8 ? _M0_0_in_waddr_T_2 : _GEN_864; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_870 = _GEN_113 == 6'h8 ? io_in_6_Im : _GEN_865; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_871 = _GEN_113 == 6'h8 ? io_in_6_Re : _GEN_866; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_874 = _GEN_130 == 6'h8 ? _M0_0_in_waddr_T_2 : _GEN_869; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_875 = _GEN_130 == 6'h8 ? io_in_7_Im : _GEN_870; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_876 = _GEN_130 == 6'h8 ? io_in_7_Re : _GEN_871; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_879 = _GEN_147 == 6'h8 ? _M0_0_in_waddr_T_26 : _GEN_874; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_880 = _GEN_147 == 6'h8 ? io_in_8_Im : _GEN_875; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_881 = _GEN_147 == 6'h8 ? io_in_8_Re : _GEN_876; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_884 = _GEN_164 == 6'h8 ? _M0_0_in_waddr_T_26 : _GEN_879; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_885 = _GEN_164 == 6'h8 ? io_in_9_Im : _GEN_880; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_886 = _GEN_164 == 6'h8 ? io_in_9_Re : _GEN_881; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_889 = _GEN_181 == 6'h8 ? _M0_0_in_waddr_T_26 : _GEN_884; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_890 = _GEN_181 == 6'h8 ? io_in_10_Im : _GEN_885; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_891 = _GEN_181 == 6'h8 ? io_in_10_Re : _GEN_886; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_894 = _GEN_198 == 6'h8 ? _M0_0_in_waddr_T_26 : _GEN_889; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_895 = _GEN_198 == 6'h8 ? io_in_11_Im : _GEN_890; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_896 = _GEN_198 == 6'h8 ? io_in_11_Re : _GEN_891; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_899 = _GEN_215 == 6'h8 ? _M0_0_in_waddr_T_26 : _GEN_894; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_900 = _GEN_215 == 6'h8 ? io_in_12_Im : _GEN_895; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_901 = _GEN_215 == 6'h8 ? io_in_12_Re : _GEN_896; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_904 = _GEN_232 == 6'h8 ? _M0_0_in_waddr_T_26 : _GEN_899; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_905 = _GEN_232 == 6'h8 ? io_in_13_Im : _GEN_900; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_906 = _GEN_232 == 6'h8 ? io_in_13_Re : _GEN_901; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_908 = _GEN_249 == 6'h8 | (_GEN_232 == 6'h8 | (_GEN_215 == 6'h8 | (_GEN_198 == 6'h8 | (_GEN_181 == 6'h8 | (
    _GEN_164 == 6'h8 | (_GEN_147 == 6'h8 | (_GEN_130 == 6'h8 | (_GEN_113 == 6'h8 | (_GEN_96 == 6'h8 | (_GEN_79 == 6'h8
     | (_GEN_62 == 6'h8 | (_GEN_45 == 6'h8 | (_GEN_28 == 6'h8 | _GEN_11 == 6'h8))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_909 = _GEN_249 == 6'h8 ? _M0_0_in_waddr_T_26 : _GEN_904; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_910 = _GEN_249 == 6'h8 ? io_in_14_Im : _GEN_905; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_911 = _GEN_249 == 6'h8 ? io_in_14_Re : _GEN_906; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_913 = _GEN_266 == 6'h8 | _GEN_908; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_914 = _GEN_266 == 6'h8 ? _M0_0_in_waddr_T_26 : _GEN_909; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_915 = _GEN_266 == 6'h8 ? io_in_15_Im : _GEN_910; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_916 = _GEN_266 == 6'h8 ? io_in_15_Re : _GEN_911; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_919 = _GEN_11 == 6'h9 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_920 = _GEN_11 == 6'h9 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_921 = _GEN_11 == 6'h9 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_924 = _GEN_28 == 6'h9 ? _M0_0_in_waddr_T_2 : _GEN_919; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_925 = _GEN_28 == 6'h9 ? io_in_1_Im : _GEN_920; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_926 = _GEN_28 == 6'h9 ? io_in_1_Re : _GEN_921; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_929 = _GEN_45 == 6'h9 ? _M0_0_in_waddr_T_2 : _GEN_924; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_930 = _GEN_45 == 6'h9 ? io_in_2_Im : _GEN_925; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_931 = _GEN_45 == 6'h9 ? io_in_2_Re : _GEN_926; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_934 = _GEN_62 == 6'h9 ? _M0_0_in_waddr_T_2 : _GEN_929; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_935 = _GEN_62 == 6'h9 ? io_in_3_Im : _GEN_930; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_936 = _GEN_62 == 6'h9 ? io_in_3_Re : _GEN_931; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_939 = _GEN_79 == 6'h9 ? _M0_0_in_waddr_T_2 : _GEN_934; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_940 = _GEN_79 == 6'h9 ? io_in_4_Im : _GEN_935; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_941 = _GEN_79 == 6'h9 ? io_in_4_Re : _GEN_936; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_944 = _GEN_96 == 6'h9 ? _M0_0_in_waddr_T_2 : _GEN_939; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_945 = _GEN_96 == 6'h9 ? io_in_5_Im : _GEN_940; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_946 = _GEN_96 == 6'h9 ? io_in_5_Re : _GEN_941; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_949 = _GEN_113 == 6'h9 ? _M0_0_in_waddr_T_2 : _GEN_944; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_950 = _GEN_113 == 6'h9 ? io_in_6_Im : _GEN_945; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_951 = _GEN_113 == 6'h9 ? io_in_6_Re : _GEN_946; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_954 = _GEN_130 == 6'h9 ? _M0_0_in_waddr_T_2 : _GEN_949; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_955 = _GEN_130 == 6'h9 ? io_in_7_Im : _GEN_950; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_956 = _GEN_130 == 6'h9 ? io_in_7_Re : _GEN_951; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_959 = _GEN_147 == 6'h9 ? _M0_0_in_waddr_T_26 : _GEN_954; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_960 = _GEN_147 == 6'h9 ? io_in_8_Im : _GEN_955; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_961 = _GEN_147 == 6'h9 ? io_in_8_Re : _GEN_956; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_964 = _GEN_164 == 6'h9 ? _M0_0_in_waddr_T_26 : _GEN_959; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_965 = _GEN_164 == 6'h9 ? io_in_9_Im : _GEN_960; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_966 = _GEN_164 == 6'h9 ? io_in_9_Re : _GEN_961; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_969 = _GEN_181 == 6'h9 ? _M0_0_in_waddr_T_26 : _GEN_964; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_970 = _GEN_181 == 6'h9 ? io_in_10_Im : _GEN_965; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_971 = _GEN_181 == 6'h9 ? io_in_10_Re : _GEN_966; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_974 = _GEN_198 == 6'h9 ? _M0_0_in_waddr_T_26 : _GEN_969; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_975 = _GEN_198 == 6'h9 ? io_in_11_Im : _GEN_970; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_976 = _GEN_198 == 6'h9 ? io_in_11_Re : _GEN_971; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_979 = _GEN_215 == 6'h9 ? _M0_0_in_waddr_T_26 : _GEN_974; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_980 = _GEN_215 == 6'h9 ? io_in_12_Im : _GEN_975; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_981 = _GEN_215 == 6'h9 ? io_in_12_Re : _GEN_976; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_984 = _GEN_232 == 6'h9 ? _M0_0_in_waddr_T_26 : _GEN_979; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_985 = _GEN_232 == 6'h9 ? io_in_13_Im : _GEN_980; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_986 = _GEN_232 == 6'h9 ? io_in_13_Re : _GEN_981; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_988 = _GEN_249 == 6'h9 | (_GEN_232 == 6'h9 | (_GEN_215 == 6'h9 | (_GEN_198 == 6'h9 | (_GEN_181 == 6'h9 | (
    _GEN_164 == 6'h9 | (_GEN_147 == 6'h9 | (_GEN_130 == 6'h9 | (_GEN_113 == 6'h9 | (_GEN_96 == 6'h9 | (_GEN_79 == 6'h9
     | (_GEN_62 == 6'h9 | (_GEN_45 == 6'h9 | (_GEN_28 == 6'h9 | _GEN_11 == 6'h9))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_989 = _GEN_249 == 6'h9 ? _M0_0_in_waddr_T_26 : _GEN_984; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_990 = _GEN_249 == 6'h9 ? io_in_14_Im : _GEN_985; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_991 = _GEN_249 == 6'h9 ? io_in_14_Re : _GEN_986; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_993 = _GEN_266 == 6'h9 | _GEN_988; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_994 = _GEN_266 == 6'h9 ? _M0_0_in_waddr_T_26 : _GEN_989; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_995 = _GEN_266 == 6'h9 ? io_in_15_Im : _GEN_990; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_996 = _GEN_266 == 6'h9 ? io_in_15_Re : _GEN_991; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_999 = _GEN_11 == 6'ha ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1000 = _GEN_11 == 6'ha ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1001 = _GEN_11 == 6'ha ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1004 = _GEN_28 == 6'ha ? _M0_0_in_waddr_T_2 : _GEN_999; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1005 = _GEN_28 == 6'ha ? io_in_1_Im : _GEN_1000; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1006 = _GEN_28 == 6'ha ? io_in_1_Re : _GEN_1001; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1009 = _GEN_45 == 6'ha ? _M0_0_in_waddr_T_2 : _GEN_1004; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1010 = _GEN_45 == 6'ha ? io_in_2_Im : _GEN_1005; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1011 = _GEN_45 == 6'ha ? io_in_2_Re : _GEN_1006; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1014 = _GEN_62 == 6'ha ? _M0_0_in_waddr_T_2 : _GEN_1009; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1015 = _GEN_62 == 6'ha ? io_in_3_Im : _GEN_1010; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1016 = _GEN_62 == 6'ha ? io_in_3_Re : _GEN_1011; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1019 = _GEN_79 == 6'ha ? _M0_0_in_waddr_T_2 : _GEN_1014; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1020 = _GEN_79 == 6'ha ? io_in_4_Im : _GEN_1015; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1021 = _GEN_79 == 6'ha ? io_in_4_Re : _GEN_1016; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1024 = _GEN_96 == 6'ha ? _M0_0_in_waddr_T_2 : _GEN_1019; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1025 = _GEN_96 == 6'ha ? io_in_5_Im : _GEN_1020; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1026 = _GEN_96 == 6'ha ? io_in_5_Re : _GEN_1021; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1029 = _GEN_113 == 6'ha ? _M0_0_in_waddr_T_2 : _GEN_1024; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1030 = _GEN_113 == 6'ha ? io_in_6_Im : _GEN_1025; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1031 = _GEN_113 == 6'ha ? io_in_6_Re : _GEN_1026; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1034 = _GEN_130 == 6'ha ? _M0_0_in_waddr_T_2 : _GEN_1029; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1035 = _GEN_130 == 6'ha ? io_in_7_Im : _GEN_1030; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1036 = _GEN_130 == 6'ha ? io_in_7_Re : _GEN_1031; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1039 = _GEN_147 == 6'ha ? _M0_0_in_waddr_T_26 : _GEN_1034; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1040 = _GEN_147 == 6'ha ? io_in_8_Im : _GEN_1035; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1041 = _GEN_147 == 6'ha ? io_in_8_Re : _GEN_1036; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1044 = _GEN_164 == 6'ha ? _M0_0_in_waddr_T_26 : _GEN_1039; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1045 = _GEN_164 == 6'ha ? io_in_9_Im : _GEN_1040; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1046 = _GEN_164 == 6'ha ? io_in_9_Re : _GEN_1041; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1049 = _GEN_181 == 6'ha ? _M0_0_in_waddr_T_26 : _GEN_1044; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1050 = _GEN_181 == 6'ha ? io_in_10_Im : _GEN_1045; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1051 = _GEN_181 == 6'ha ? io_in_10_Re : _GEN_1046; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1054 = _GEN_198 == 6'ha ? _M0_0_in_waddr_T_26 : _GEN_1049; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1055 = _GEN_198 == 6'ha ? io_in_11_Im : _GEN_1050; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1056 = _GEN_198 == 6'ha ? io_in_11_Re : _GEN_1051; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1059 = _GEN_215 == 6'ha ? _M0_0_in_waddr_T_26 : _GEN_1054; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1060 = _GEN_215 == 6'ha ? io_in_12_Im : _GEN_1055; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1061 = _GEN_215 == 6'ha ? io_in_12_Re : _GEN_1056; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1064 = _GEN_232 == 6'ha ? _M0_0_in_waddr_T_26 : _GEN_1059; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1065 = _GEN_232 == 6'ha ? io_in_13_Im : _GEN_1060; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1066 = _GEN_232 == 6'ha ? io_in_13_Re : _GEN_1061; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1068 = _GEN_249 == 6'ha | (_GEN_232 == 6'ha | (_GEN_215 == 6'ha | (_GEN_198 == 6'ha | (_GEN_181 == 6'ha | (
    _GEN_164 == 6'ha | (_GEN_147 == 6'ha | (_GEN_130 == 6'ha | (_GEN_113 == 6'ha | (_GEN_96 == 6'ha | (_GEN_79 == 6'ha
     | (_GEN_62 == 6'ha | (_GEN_45 == 6'ha | (_GEN_28 == 6'ha | _GEN_11 == 6'ha))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1069 = _GEN_249 == 6'ha ? _M0_0_in_waddr_T_26 : _GEN_1064; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1070 = _GEN_249 == 6'ha ? io_in_14_Im : _GEN_1065; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1071 = _GEN_249 == 6'ha ? io_in_14_Re : _GEN_1066; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1073 = _GEN_266 == 6'ha | _GEN_1068; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1074 = _GEN_266 == 6'ha ? _M0_0_in_waddr_T_26 : _GEN_1069; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1075 = _GEN_266 == 6'ha ? io_in_15_Im : _GEN_1070; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1076 = _GEN_266 == 6'ha ? io_in_15_Re : _GEN_1071; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1079 = _GEN_11 == 6'hb ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1080 = _GEN_11 == 6'hb ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1081 = _GEN_11 == 6'hb ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1084 = _GEN_28 == 6'hb ? _M0_0_in_waddr_T_2 : _GEN_1079; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1085 = _GEN_28 == 6'hb ? io_in_1_Im : _GEN_1080; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1086 = _GEN_28 == 6'hb ? io_in_1_Re : _GEN_1081; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1089 = _GEN_45 == 6'hb ? _M0_0_in_waddr_T_2 : _GEN_1084; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1090 = _GEN_45 == 6'hb ? io_in_2_Im : _GEN_1085; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1091 = _GEN_45 == 6'hb ? io_in_2_Re : _GEN_1086; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1094 = _GEN_62 == 6'hb ? _M0_0_in_waddr_T_2 : _GEN_1089; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1095 = _GEN_62 == 6'hb ? io_in_3_Im : _GEN_1090; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1096 = _GEN_62 == 6'hb ? io_in_3_Re : _GEN_1091; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1099 = _GEN_79 == 6'hb ? _M0_0_in_waddr_T_2 : _GEN_1094; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1100 = _GEN_79 == 6'hb ? io_in_4_Im : _GEN_1095; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1101 = _GEN_79 == 6'hb ? io_in_4_Re : _GEN_1096; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1104 = _GEN_96 == 6'hb ? _M0_0_in_waddr_T_2 : _GEN_1099; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1105 = _GEN_96 == 6'hb ? io_in_5_Im : _GEN_1100; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1106 = _GEN_96 == 6'hb ? io_in_5_Re : _GEN_1101; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1109 = _GEN_113 == 6'hb ? _M0_0_in_waddr_T_2 : _GEN_1104; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1110 = _GEN_113 == 6'hb ? io_in_6_Im : _GEN_1105; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1111 = _GEN_113 == 6'hb ? io_in_6_Re : _GEN_1106; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1114 = _GEN_130 == 6'hb ? _M0_0_in_waddr_T_2 : _GEN_1109; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1115 = _GEN_130 == 6'hb ? io_in_7_Im : _GEN_1110; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1116 = _GEN_130 == 6'hb ? io_in_7_Re : _GEN_1111; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1119 = _GEN_147 == 6'hb ? _M0_0_in_waddr_T_26 : _GEN_1114; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1120 = _GEN_147 == 6'hb ? io_in_8_Im : _GEN_1115; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1121 = _GEN_147 == 6'hb ? io_in_8_Re : _GEN_1116; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1124 = _GEN_164 == 6'hb ? _M0_0_in_waddr_T_26 : _GEN_1119; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1125 = _GEN_164 == 6'hb ? io_in_9_Im : _GEN_1120; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1126 = _GEN_164 == 6'hb ? io_in_9_Re : _GEN_1121; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1129 = _GEN_181 == 6'hb ? _M0_0_in_waddr_T_26 : _GEN_1124; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1130 = _GEN_181 == 6'hb ? io_in_10_Im : _GEN_1125; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1131 = _GEN_181 == 6'hb ? io_in_10_Re : _GEN_1126; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1134 = _GEN_198 == 6'hb ? _M0_0_in_waddr_T_26 : _GEN_1129; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1135 = _GEN_198 == 6'hb ? io_in_11_Im : _GEN_1130; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1136 = _GEN_198 == 6'hb ? io_in_11_Re : _GEN_1131; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1139 = _GEN_215 == 6'hb ? _M0_0_in_waddr_T_26 : _GEN_1134; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1140 = _GEN_215 == 6'hb ? io_in_12_Im : _GEN_1135; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1141 = _GEN_215 == 6'hb ? io_in_12_Re : _GEN_1136; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1144 = _GEN_232 == 6'hb ? _M0_0_in_waddr_T_26 : _GEN_1139; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1145 = _GEN_232 == 6'hb ? io_in_13_Im : _GEN_1140; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1146 = _GEN_232 == 6'hb ? io_in_13_Re : _GEN_1141; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1148 = _GEN_249 == 6'hb | (_GEN_232 == 6'hb | (_GEN_215 == 6'hb | (_GEN_198 == 6'hb | (_GEN_181 == 6'hb | (
    _GEN_164 == 6'hb | (_GEN_147 == 6'hb | (_GEN_130 == 6'hb | (_GEN_113 == 6'hb | (_GEN_96 == 6'hb | (_GEN_79 == 6'hb
     | (_GEN_62 == 6'hb | (_GEN_45 == 6'hb | (_GEN_28 == 6'hb | _GEN_11 == 6'hb))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1149 = _GEN_249 == 6'hb ? _M0_0_in_waddr_T_26 : _GEN_1144; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1150 = _GEN_249 == 6'hb ? io_in_14_Im : _GEN_1145; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1151 = _GEN_249 == 6'hb ? io_in_14_Re : _GEN_1146; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1153 = _GEN_266 == 6'hb | _GEN_1148; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1154 = _GEN_266 == 6'hb ? _M0_0_in_waddr_T_26 : _GEN_1149; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1155 = _GEN_266 == 6'hb ? io_in_15_Im : _GEN_1150; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1156 = _GEN_266 == 6'hb ? io_in_15_Re : _GEN_1151; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1159 = _GEN_11 == 6'hc ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1160 = _GEN_11 == 6'hc ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1161 = _GEN_11 == 6'hc ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1164 = _GEN_28 == 6'hc ? _M0_0_in_waddr_T_2 : _GEN_1159; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1165 = _GEN_28 == 6'hc ? io_in_1_Im : _GEN_1160; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1166 = _GEN_28 == 6'hc ? io_in_1_Re : _GEN_1161; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1169 = _GEN_45 == 6'hc ? _M0_0_in_waddr_T_2 : _GEN_1164; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1170 = _GEN_45 == 6'hc ? io_in_2_Im : _GEN_1165; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1171 = _GEN_45 == 6'hc ? io_in_2_Re : _GEN_1166; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1174 = _GEN_62 == 6'hc ? _M0_0_in_waddr_T_2 : _GEN_1169; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1175 = _GEN_62 == 6'hc ? io_in_3_Im : _GEN_1170; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1176 = _GEN_62 == 6'hc ? io_in_3_Re : _GEN_1171; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1179 = _GEN_79 == 6'hc ? _M0_0_in_waddr_T_2 : _GEN_1174; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1180 = _GEN_79 == 6'hc ? io_in_4_Im : _GEN_1175; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1181 = _GEN_79 == 6'hc ? io_in_4_Re : _GEN_1176; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1184 = _GEN_96 == 6'hc ? _M0_0_in_waddr_T_2 : _GEN_1179; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1185 = _GEN_96 == 6'hc ? io_in_5_Im : _GEN_1180; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1186 = _GEN_96 == 6'hc ? io_in_5_Re : _GEN_1181; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1189 = _GEN_113 == 6'hc ? _M0_0_in_waddr_T_2 : _GEN_1184; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1190 = _GEN_113 == 6'hc ? io_in_6_Im : _GEN_1185; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1191 = _GEN_113 == 6'hc ? io_in_6_Re : _GEN_1186; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1194 = _GEN_130 == 6'hc ? _M0_0_in_waddr_T_2 : _GEN_1189; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1195 = _GEN_130 == 6'hc ? io_in_7_Im : _GEN_1190; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1196 = _GEN_130 == 6'hc ? io_in_7_Re : _GEN_1191; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1199 = _GEN_147 == 6'hc ? _M0_0_in_waddr_T_26 : _GEN_1194; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1200 = _GEN_147 == 6'hc ? io_in_8_Im : _GEN_1195; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1201 = _GEN_147 == 6'hc ? io_in_8_Re : _GEN_1196; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1204 = _GEN_164 == 6'hc ? _M0_0_in_waddr_T_26 : _GEN_1199; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1205 = _GEN_164 == 6'hc ? io_in_9_Im : _GEN_1200; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1206 = _GEN_164 == 6'hc ? io_in_9_Re : _GEN_1201; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1209 = _GEN_181 == 6'hc ? _M0_0_in_waddr_T_26 : _GEN_1204; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1210 = _GEN_181 == 6'hc ? io_in_10_Im : _GEN_1205; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1211 = _GEN_181 == 6'hc ? io_in_10_Re : _GEN_1206; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1214 = _GEN_198 == 6'hc ? _M0_0_in_waddr_T_26 : _GEN_1209; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1215 = _GEN_198 == 6'hc ? io_in_11_Im : _GEN_1210; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1216 = _GEN_198 == 6'hc ? io_in_11_Re : _GEN_1211; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1219 = _GEN_215 == 6'hc ? _M0_0_in_waddr_T_26 : _GEN_1214; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1220 = _GEN_215 == 6'hc ? io_in_12_Im : _GEN_1215; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1221 = _GEN_215 == 6'hc ? io_in_12_Re : _GEN_1216; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1224 = _GEN_232 == 6'hc ? _M0_0_in_waddr_T_26 : _GEN_1219; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1225 = _GEN_232 == 6'hc ? io_in_13_Im : _GEN_1220; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1226 = _GEN_232 == 6'hc ? io_in_13_Re : _GEN_1221; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1228 = _GEN_249 == 6'hc | (_GEN_232 == 6'hc | (_GEN_215 == 6'hc | (_GEN_198 == 6'hc | (_GEN_181 == 6'hc | (
    _GEN_164 == 6'hc | (_GEN_147 == 6'hc | (_GEN_130 == 6'hc | (_GEN_113 == 6'hc | (_GEN_96 == 6'hc | (_GEN_79 == 6'hc
     | (_GEN_62 == 6'hc | (_GEN_45 == 6'hc | (_GEN_28 == 6'hc | _GEN_11 == 6'hc))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1229 = _GEN_249 == 6'hc ? _M0_0_in_waddr_T_26 : _GEN_1224; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1230 = _GEN_249 == 6'hc ? io_in_14_Im : _GEN_1225; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1231 = _GEN_249 == 6'hc ? io_in_14_Re : _GEN_1226; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1233 = _GEN_266 == 6'hc | _GEN_1228; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1234 = _GEN_266 == 6'hc ? _M0_0_in_waddr_T_26 : _GEN_1229; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1235 = _GEN_266 == 6'hc ? io_in_15_Im : _GEN_1230; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1236 = _GEN_266 == 6'hc ? io_in_15_Re : _GEN_1231; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1239 = _GEN_11 == 6'hd ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1240 = _GEN_11 == 6'hd ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1241 = _GEN_11 == 6'hd ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1244 = _GEN_28 == 6'hd ? _M0_0_in_waddr_T_2 : _GEN_1239; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1245 = _GEN_28 == 6'hd ? io_in_1_Im : _GEN_1240; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1246 = _GEN_28 == 6'hd ? io_in_1_Re : _GEN_1241; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1249 = _GEN_45 == 6'hd ? _M0_0_in_waddr_T_2 : _GEN_1244; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1250 = _GEN_45 == 6'hd ? io_in_2_Im : _GEN_1245; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1251 = _GEN_45 == 6'hd ? io_in_2_Re : _GEN_1246; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1254 = _GEN_62 == 6'hd ? _M0_0_in_waddr_T_2 : _GEN_1249; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1255 = _GEN_62 == 6'hd ? io_in_3_Im : _GEN_1250; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1256 = _GEN_62 == 6'hd ? io_in_3_Re : _GEN_1251; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1259 = _GEN_79 == 6'hd ? _M0_0_in_waddr_T_2 : _GEN_1254; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1260 = _GEN_79 == 6'hd ? io_in_4_Im : _GEN_1255; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1261 = _GEN_79 == 6'hd ? io_in_4_Re : _GEN_1256; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1264 = _GEN_96 == 6'hd ? _M0_0_in_waddr_T_2 : _GEN_1259; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1265 = _GEN_96 == 6'hd ? io_in_5_Im : _GEN_1260; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1266 = _GEN_96 == 6'hd ? io_in_5_Re : _GEN_1261; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1269 = _GEN_113 == 6'hd ? _M0_0_in_waddr_T_2 : _GEN_1264; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1270 = _GEN_113 == 6'hd ? io_in_6_Im : _GEN_1265; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1271 = _GEN_113 == 6'hd ? io_in_6_Re : _GEN_1266; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1274 = _GEN_130 == 6'hd ? _M0_0_in_waddr_T_2 : _GEN_1269; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1275 = _GEN_130 == 6'hd ? io_in_7_Im : _GEN_1270; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1276 = _GEN_130 == 6'hd ? io_in_7_Re : _GEN_1271; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1279 = _GEN_147 == 6'hd ? _M0_0_in_waddr_T_26 : _GEN_1274; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1280 = _GEN_147 == 6'hd ? io_in_8_Im : _GEN_1275; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1281 = _GEN_147 == 6'hd ? io_in_8_Re : _GEN_1276; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1284 = _GEN_164 == 6'hd ? _M0_0_in_waddr_T_26 : _GEN_1279; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1285 = _GEN_164 == 6'hd ? io_in_9_Im : _GEN_1280; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1286 = _GEN_164 == 6'hd ? io_in_9_Re : _GEN_1281; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1289 = _GEN_181 == 6'hd ? _M0_0_in_waddr_T_26 : _GEN_1284; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1290 = _GEN_181 == 6'hd ? io_in_10_Im : _GEN_1285; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1291 = _GEN_181 == 6'hd ? io_in_10_Re : _GEN_1286; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1294 = _GEN_198 == 6'hd ? _M0_0_in_waddr_T_26 : _GEN_1289; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1295 = _GEN_198 == 6'hd ? io_in_11_Im : _GEN_1290; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1296 = _GEN_198 == 6'hd ? io_in_11_Re : _GEN_1291; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1299 = _GEN_215 == 6'hd ? _M0_0_in_waddr_T_26 : _GEN_1294; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1300 = _GEN_215 == 6'hd ? io_in_12_Im : _GEN_1295; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1301 = _GEN_215 == 6'hd ? io_in_12_Re : _GEN_1296; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1304 = _GEN_232 == 6'hd ? _M0_0_in_waddr_T_26 : _GEN_1299; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1305 = _GEN_232 == 6'hd ? io_in_13_Im : _GEN_1300; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1306 = _GEN_232 == 6'hd ? io_in_13_Re : _GEN_1301; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1308 = _GEN_249 == 6'hd | (_GEN_232 == 6'hd | (_GEN_215 == 6'hd | (_GEN_198 == 6'hd | (_GEN_181 == 6'hd | (
    _GEN_164 == 6'hd | (_GEN_147 == 6'hd | (_GEN_130 == 6'hd | (_GEN_113 == 6'hd | (_GEN_96 == 6'hd | (_GEN_79 == 6'hd
     | (_GEN_62 == 6'hd | (_GEN_45 == 6'hd | (_GEN_28 == 6'hd | _GEN_11 == 6'hd))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1309 = _GEN_249 == 6'hd ? _M0_0_in_waddr_T_26 : _GEN_1304; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1310 = _GEN_249 == 6'hd ? io_in_14_Im : _GEN_1305; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1311 = _GEN_249 == 6'hd ? io_in_14_Re : _GEN_1306; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1313 = _GEN_266 == 6'hd | _GEN_1308; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1314 = _GEN_266 == 6'hd ? _M0_0_in_waddr_T_26 : _GEN_1309; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1315 = _GEN_266 == 6'hd ? io_in_15_Im : _GEN_1310; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1316 = _GEN_266 == 6'hd ? io_in_15_Re : _GEN_1311; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1319 = _GEN_11 == 6'he ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1320 = _GEN_11 == 6'he ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1321 = _GEN_11 == 6'he ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1324 = _GEN_28 == 6'he ? _M0_0_in_waddr_T_2 : _GEN_1319; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1325 = _GEN_28 == 6'he ? io_in_1_Im : _GEN_1320; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1326 = _GEN_28 == 6'he ? io_in_1_Re : _GEN_1321; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1329 = _GEN_45 == 6'he ? _M0_0_in_waddr_T_2 : _GEN_1324; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1330 = _GEN_45 == 6'he ? io_in_2_Im : _GEN_1325; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1331 = _GEN_45 == 6'he ? io_in_2_Re : _GEN_1326; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1334 = _GEN_62 == 6'he ? _M0_0_in_waddr_T_2 : _GEN_1329; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1335 = _GEN_62 == 6'he ? io_in_3_Im : _GEN_1330; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1336 = _GEN_62 == 6'he ? io_in_3_Re : _GEN_1331; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1339 = _GEN_79 == 6'he ? _M0_0_in_waddr_T_2 : _GEN_1334; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1340 = _GEN_79 == 6'he ? io_in_4_Im : _GEN_1335; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1341 = _GEN_79 == 6'he ? io_in_4_Re : _GEN_1336; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1344 = _GEN_96 == 6'he ? _M0_0_in_waddr_T_2 : _GEN_1339; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1345 = _GEN_96 == 6'he ? io_in_5_Im : _GEN_1340; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1346 = _GEN_96 == 6'he ? io_in_5_Re : _GEN_1341; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1349 = _GEN_113 == 6'he ? _M0_0_in_waddr_T_2 : _GEN_1344; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1350 = _GEN_113 == 6'he ? io_in_6_Im : _GEN_1345; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1351 = _GEN_113 == 6'he ? io_in_6_Re : _GEN_1346; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1354 = _GEN_130 == 6'he ? _M0_0_in_waddr_T_2 : _GEN_1349; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1355 = _GEN_130 == 6'he ? io_in_7_Im : _GEN_1350; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1356 = _GEN_130 == 6'he ? io_in_7_Re : _GEN_1351; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1359 = _GEN_147 == 6'he ? _M0_0_in_waddr_T_26 : _GEN_1354; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1360 = _GEN_147 == 6'he ? io_in_8_Im : _GEN_1355; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1361 = _GEN_147 == 6'he ? io_in_8_Re : _GEN_1356; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1364 = _GEN_164 == 6'he ? _M0_0_in_waddr_T_26 : _GEN_1359; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1365 = _GEN_164 == 6'he ? io_in_9_Im : _GEN_1360; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1366 = _GEN_164 == 6'he ? io_in_9_Re : _GEN_1361; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1369 = _GEN_181 == 6'he ? _M0_0_in_waddr_T_26 : _GEN_1364; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1370 = _GEN_181 == 6'he ? io_in_10_Im : _GEN_1365; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1371 = _GEN_181 == 6'he ? io_in_10_Re : _GEN_1366; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1374 = _GEN_198 == 6'he ? _M0_0_in_waddr_T_26 : _GEN_1369; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1375 = _GEN_198 == 6'he ? io_in_11_Im : _GEN_1370; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1376 = _GEN_198 == 6'he ? io_in_11_Re : _GEN_1371; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1379 = _GEN_215 == 6'he ? _M0_0_in_waddr_T_26 : _GEN_1374; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1380 = _GEN_215 == 6'he ? io_in_12_Im : _GEN_1375; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1381 = _GEN_215 == 6'he ? io_in_12_Re : _GEN_1376; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1384 = _GEN_232 == 6'he ? _M0_0_in_waddr_T_26 : _GEN_1379; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1385 = _GEN_232 == 6'he ? io_in_13_Im : _GEN_1380; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1386 = _GEN_232 == 6'he ? io_in_13_Re : _GEN_1381; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1388 = _GEN_249 == 6'he | (_GEN_232 == 6'he | (_GEN_215 == 6'he | (_GEN_198 == 6'he | (_GEN_181 == 6'he | (
    _GEN_164 == 6'he | (_GEN_147 == 6'he | (_GEN_130 == 6'he | (_GEN_113 == 6'he | (_GEN_96 == 6'he | (_GEN_79 == 6'he
     | (_GEN_62 == 6'he | (_GEN_45 == 6'he | (_GEN_28 == 6'he | _GEN_11 == 6'he))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1389 = _GEN_249 == 6'he ? _M0_0_in_waddr_T_26 : _GEN_1384; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1390 = _GEN_249 == 6'he ? io_in_14_Im : _GEN_1385; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1391 = _GEN_249 == 6'he ? io_in_14_Re : _GEN_1386; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1393 = _GEN_266 == 6'he | _GEN_1388; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1394 = _GEN_266 == 6'he ? _M0_0_in_waddr_T_26 : _GEN_1389; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1395 = _GEN_266 == 6'he ? io_in_15_Im : _GEN_1390; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1396 = _GEN_266 == 6'he ? io_in_15_Re : _GEN_1391; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1399 = _GEN_11 == 6'hf ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1400 = _GEN_11 == 6'hf ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1401 = _GEN_11 == 6'hf ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1404 = _GEN_28 == 6'hf ? _M0_0_in_waddr_T_2 : _GEN_1399; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1405 = _GEN_28 == 6'hf ? io_in_1_Im : _GEN_1400; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1406 = _GEN_28 == 6'hf ? io_in_1_Re : _GEN_1401; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1409 = _GEN_45 == 6'hf ? _M0_0_in_waddr_T_2 : _GEN_1404; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1410 = _GEN_45 == 6'hf ? io_in_2_Im : _GEN_1405; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1411 = _GEN_45 == 6'hf ? io_in_2_Re : _GEN_1406; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1414 = _GEN_62 == 6'hf ? _M0_0_in_waddr_T_2 : _GEN_1409; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1415 = _GEN_62 == 6'hf ? io_in_3_Im : _GEN_1410; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1416 = _GEN_62 == 6'hf ? io_in_3_Re : _GEN_1411; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1419 = _GEN_79 == 6'hf ? _M0_0_in_waddr_T_2 : _GEN_1414; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1420 = _GEN_79 == 6'hf ? io_in_4_Im : _GEN_1415; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1421 = _GEN_79 == 6'hf ? io_in_4_Re : _GEN_1416; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1424 = _GEN_96 == 6'hf ? _M0_0_in_waddr_T_2 : _GEN_1419; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1425 = _GEN_96 == 6'hf ? io_in_5_Im : _GEN_1420; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1426 = _GEN_96 == 6'hf ? io_in_5_Re : _GEN_1421; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1429 = _GEN_113 == 6'hf ? _M0_0_in_waddr_T_2 : _GEN_1424; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1430 = _GEN_113 == 6'hf ? io_in_6_Im : _GEN_1425; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1431 = _GEN_113 == 6'hf ? io_in_6_Re : _GEN_1426; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1434 = _GEN_130 == 6'hf ? _M0_0_in_waddr_T_2 : _GEN_1429; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1435 = _GEN_130 == 6'hf ? io_in_7_Im : _GEN_1430; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1436 = _GEN_130 == 6'hf ? io_in_7_Re : _GEN_1431; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1439 = _GEN_147 == 6'hf ? _M0_0_in_waddr_T_26 : _GEN_1434; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1440 = _GEN_147 == 6'hf ? io_in_8_Im : _GEN_1435; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1441 = _GEN_147 == 6'hf ? io_in_8_Re : _GEN_1436; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1444 = _GEN_164 == 6'hf ? _M0_0_in_waddr_T_26 : _GEN_1439; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1445 = _GEN_164 == 6'hf ? io_in_9_Im : _GEN_1440; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1446 = _GEN_164 == 6'hf ? io_in_9_Re : _GEN_1441; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1449 = _GEN_181 == 6'hf ? _M0_0_in_waddr_T_26 : _GEN_1444; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1450 = _GEN_181 == 6'hf ? io_in_10_Im : _GEN_1445; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1451 = _GEN_181 == 6'hf ? io_in_10_Re : _GEN_1446; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1454 = _GEN_198 == 6'hf ? _M0_0_in_waddr_T_26 : _GEN_1449; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1455 = _GEN_198 == 6'hf ? io_in_11_Im : _GEN_1450; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1456 = _GEN_198 == 6'hf ? io_in_11_Re : _GEN_1451; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1459 = _GEN_215 == 6'hf ? _M0_0_in_waddr_T_26 : _GEN_1454; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1460 = _GEN_215 == 6'hf ? io_in_12_Im : _GEN_1455; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1461 = _GEN_215 == 6'hf ? io_in_12_Re : _GEN_1456; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1464 = _GEN_232 == 6'hf ? _M0_0_in_waddr_T_26 : _GEN_1459; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1465 = _GEN_232 == 6'hf ? io_in_13_Im : _GEN_1460; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1466 = _GEN_232 == 6'hf ? io_in_13_Re : _GEN_1461; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1468 = _GEN_249 == 6'hf | (_GEN_232 == 6'hf | (_GEN_215 == 6'hf | (_GEN_198 == 6'hf | (_GEN_181 == 6'hf | (
    _GEN_164 == 6'hf | (_GEN_147 == 6'hf | (_GEN_130 == 6'hf | (_GEN_113 == 6'hf | (_GEN_96 == 6'hf | (_GEN_79 == 6'hf
     | (_GEN_62 == 6'hf | (_GEN_45 == 6'hf | (_GEN_28 == 6'hf | _GEN_11 == 6'hf))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1469 = _GEN_249 == 6'hf ? _M0_0_in_waddr_T_26 : _GEN_1464; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1470 = _GEN_249 == 6'hf ? io_in_14_Im : _GEN_1465; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1471 = _GEN_249 == 6'hf ? io_in_14_Re : _GEN_1466; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1473 = _GEN_266 == 6'hf | _GEN_1468; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1474 = _GEN_266 == 6'hf ? _M0_0_in_waddr_T_26 : _GEN_1469; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1475 = _GEN_266 == 6'hf ? io_in_15_Im : _GEN_1470; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1476 = _GEN_266 == 6'hf ? io_in_15_Re : _GEN_1471; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1479 = _GEN_11 == 6'h10 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1480 = _GEN_11 == 6'h10 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1481 = _GEN_11 == 6'h10 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1484 = _GEN_28 == 6'h10 ? _M0_0_in_waddr_T_2 : _GEN_1479; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1485 = _GEN_28 == 6'h10 ? io_in_1_Im : _GEN_1480; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1486 = _GEN_28 == 6'h10 ? io_in_1_Re : _GEN_1481; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1489 = _GEN_45 == 6'h10 ? _M0_0_in_waddr_T_2 : _GEN_1484; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1490 = _GEN_45 == 6'h10 ? io_in_2_Im : _GEN_1485; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1491 = _GEN_45 == 6'h10 ? io_in_2_Re : _GEN_1486; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1494 = _GEN_62 == 6'h10 ? _M0_0_in_waddr_T_2 : _GEN_1489; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1495 = _GEN_62 == 6'h10 ? io_in_3_Im : _GEN_1490; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1496 = _GEN_62 == 6'h10 ? io_in_3_Re : _GEN_1491; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1499 = _GEN_79 == 6'h10 ? _M0_0_in_waddr_T_2 : _GEN_1494; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1500 = _GEN_79 == 6'h10 ? io_in_4_Im : _GEN_1495; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1501 = _GEN_79 == 6'h10 ? io_in_4_Re : _GEN_1496; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1504 = _GEN_96 == 6'h10 ? _M0_0_in_waddr_T_2 : _GEN_1499; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1505 = _GEN_96 == 6'h10 ? io_in_5_Im : _GEN_1500; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1506 = _GEN_96 == 6'h10 ? io_in_5_Re : _GEN_1501; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1509 = _GEN_113 == 6'h10 ? _M0_0_in_waddr_T_2 : _GEN_1504; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1510 = _GEN_113 == 6'h10 ? io_in_6_Im : _GEN_1505; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1511 = _GEN_113 == 6'h10 ? io_in_6_Re : _GEN_1506; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1514 = _GEN_130 == 6'h10 ? _M0_0_in_waddr_T_2 : _GEN_1509; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1515 = _GEN_130 == 6'h10 ? io_in_7_Im : _GEN_1510; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1516 = _GEN_130 == 6'h10 ? io_in_7_Re : _GEN_1511; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1519 = _GEN_147 == 6'h10 ? _M0_0_in_waddr_T_26 : _GEN_1514; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1520 = _GEN_147 == 6'h10 ? io_in_8_Im : _GEN_1515; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1521 = _GEN_147 == 6'h10 ? io_in_8_Re : _GEN_1516; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1524 = _GEN_164 == 6'h10 ? _M0_0_in_waddr_T_26 : _GEN_1519; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1525 = _GEN_164 == 6'h10 ? io_in_9_Im : _GEN_1520; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1526 = _GEN_164 == 6'h10 ? io_in_9_Re : _GEN_1521; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1529 = _GEN_181 == 6'h10 ? _M0_0_in_waddr_T_26 : _GEN_1524; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1530 = _GEN_181 == 6'h10 ? io_in_10_Im : _GEN_1525; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1531 = _GEN_181 == 6'h10 ? io_in_10_Re : _GEN_1526; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1534 = _GEN_198 == 6'h10 ? _M0_0_in_waddr_T_26 : _GEN_1529; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1535 = _GEN_198 == 6'h10 ? io_in_11_Im : _GEN_1530; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1536 = _GEN_198 == 6'h10 ? io_in_11_Re : _GEN_1531; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1539 = _GEN_215 == 6'h10 ? _M0_0_in_waddr_T_26 : _GEN_1534; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1540 = _GEN_215 == 6'h10 ? io_in_12_Im : _GEN_1535; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1541 = _GEN_215 == 6'h10 ? io_in_12_Re : _GEN_1536; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1544 = _GEN_232 == 6'h10 ? _M0_0_in_waddr_T_26 : _GEN_1539; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1545 = _GEN_232 == 6'h10 ? io_in_13_Im : _GEN_1540; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1546 = _GEN_232 == 6'h10 ? io_in_13_Re : _GEN_1541; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1548 = _GEN_249 == 6'h10 | (_GEN_232 == 6'h10 | (_GEN_215 == 6'h10 | (_GEN_198 == 6'h10 | (_GEN_181 == 6'h10
     | (_GEN_164 == 6'h10 | (_GEN_147 == 6'h10 | (_GEN_130 == 6'h10 | (_GEN_113 == 6'h10 | (_GEN_96 == 6'h10 | (_GEN_79
     == 6'h10 | (_GEN_62 == 6'h10 | (_GEN_45 == 6'h10 | (_GEN_28 == 6'h10 | _GEN_11 == 6'h10))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1549 = _GEN_249 == 6'h10 ? _M0_0_in_waddr_T_26 : _GEN_1544; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1550 = _GEN_249 == 6'h10 ? io_in_14_Im : _GEN_1545; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1551 = _GEN_249 == 6'h10 ? io_in_14_Re : _GEN_1546; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1553 = _GEN_266 == 6'h10 | _GEN_1548; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1554 = _GEN_266 == 6'h10 ? _M0_0_in_waddr_T_26 : _GEN_1549; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1555 = _GEN_266 == 6'h10 ? io_in_15_Im : _GEN_1550; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1556 = _GEN_266 == 6'h10 ? io_in_15_Re : _GEN_1551; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1559 = _GEN_11 == 6'h11 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1560 = _GEN_11 == 6'h11 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1561 = _GEN_11 == 6'h11 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1564 = _GEN_28 == 6'h11 ? _M0_0_in_waddr_T_2 : _GEN_1559; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1565 = _GEN_28 == 6'h11 ? io_in_1_Im : _GEN_1560; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1566 = _GEN_28 == 6'h11 ? io_in_1_Re : _GEN_1561; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1569 = _GEN_45 == 6'h11 ? _M0_0_in_waddr_T_2 : _GEN_1564; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1570 = _GEN_45 == 6'h11 ? io_in_2_Im : _GEN_1565; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1571 = _GEN_45 == 6'h11 ? io_in_2_Re : _GEN_1566; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1574 = _GEN_62 == 6'h11 ? _M0_0_in_waddr_T_2 : _GEN_1569; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1575 = _GEN_62 == 6'h11 ? io_in_3_Im : _GEN_1570; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1576 = _GEN_62 == 6'h11 ? io_in_3_Re : _GEN_1571; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1579 = _GEN_79 == 6'h11 ? _M0_0_in_waddr_T_2 : _GEN_1574; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1580 = _GEN_79 == 6'h11 ? io_in_4_Im : _GEN_1575; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1581 = _GEN_79 == 6'h11 ? io_in_4_Re : _GEN_1576; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1584 = _GEN_96 == 6'h11 ? _M0_0_in_waddr_T_2 : _GEN_1579; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1585 = _GEN_96 == 6'h11 ? io_in_5_Im : _GEN_1580; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1586 = _GEN_96 == 6'h11 ? io_in_5_Re : _GEN_1581; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1589 = _GEN_113 == 6'h11 ? _M0_0_in_waddr_T_2 : _GEN_1584; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1590 = _GEN_113 == 6'h11 ? io_in_6_Im : _GEN_1585; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1591 = _GEN_113 == 6'h11 ? io_in_6_Re : _GEN_1586; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1594 = _GEN_130 == 6'h11 ? _M0_0_in_waddr_T_2 : _GEN_1589; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1595 = _GEN_130 == 6'h11 ? io_in_7_Im : _GEN_1590; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1596 = _GEN_130 == 6'h11 ? io_in_7_Re : _GEN_1591; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1599 = _GEN_147 == 6'h11 ? _M0_0_in_waddr_T_26 : _GEN_1594; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1600 = _GEN_147 == 6'h11 ? io_in_8_Im : _GEN_1595; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1601 = _GEN_147 == 6'h11 ? io_in_8_Re : _GEN_1596; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1604 = _GEN_164 == 6'h11 ? _M0_0_in_waddr_T_26 : _GEN_1599; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1605 = _GEN_164 == 6'h11 ? io_in_9_Im : _GEN_1600; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1606 = _GEN_164 == 6'h11 ? io_in_9_Re : _GEN_1601; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1609 = _GEN_181 == 6'h11 ? _M0_0_in_waddr_T_26 : _GEN_1604; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1610 = _GEN_181 == 6'h11 ? io_in_10_Im : _GEN_1605; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1611 = _GEN_181 == 6'h11 ? io_in_10_Re : _GEN_1606; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1614 = _GEN_198 == 6'h11 ? _M0_0_in_waddr_T_26 : _GEN_1609; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1615 = _GEN_198 == 6'h11 ? io_in_11_Im : _GEN_1610; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1616 = _GEN_198 == 6'h11 ? io_in_11_Re : _GEN_1611; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1619 = _GEN_215 == 6'h11 ? _M0_0_in_waddr_T_26 : _GEN_1614; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1620 = _GEN_215 == 6'h11 ? io_in_12_Im : _GEN_1615; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1621 = _GEN_215 == 6'h11 ? io_in_12_Re : _GEN_1616; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1624 = _GEN_232 == 6'h11 ? _M0_0_in_waddr_T_26 : _GEN_1619; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1625 = _GEN_232 == 6'h11 ? io_in_13_Im : _GEN_1620; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1626 = _GEN_232 == 6'h11 ? io_in_13_Re : _GEN_1621; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1628 = _GEN_249 == 6'h11 | (_GEN_232 == 6'h11 | (_GEN_215 == 6'h11 | (_GEN_198 == 6'h11 | (_GEN_181 == 6'h11
     | (_GEN_164 == 6'h11 | (_GEN_147 == 6'h11 | (_GEN_130 == 6'h11 | (_GEN_113 == 6'h11 | (_GEN_96 == 6'h11 | (_GEN_79
     == 6'h11 | (_GEN_62 == 6'h11 | (_GEN_45 == 6'h11 | (_GEN_28 == 6'h11 | _GEN_11 == 6'h11))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1629 = _GEN_249 == 6'h11 ? _M0_0_in_waddr_T_26 : _GEN_1624; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1630 = _GEN_249 == 6'h11 ? io_in_14_Im : _GEN_1625; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1631 = _GEN_249 == 6'h11 ? io_in_14_Re : _GEN_1626; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1633 = _GEN_266 == 6'h11 | _GEN_1628; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1634 = _GEN_266 == 6'h11 ? _M0_0_in_waddr_T_26 : _GEN_1629; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1635 = _GEN_266 == 6'h11 ? io_in_15_Im : _GEN_1630; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1636 = _GEN_266 == 6'h11 ? io_in_15_Re : _GEN_1631; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1639 = _GEN_11 == 6'h12 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1640 = _GEN_11 == 6'h12 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1641 = _GEN_11 == 6'h12 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1644 = _GEN_28 == 6'h12 ? _M0_0_in_waddr_T_2 : _GEN_1639; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1645 = _GEN_28 == 6'h12 ? io_in_1_Im : _GEN_1640; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1646 = _GEN_28 == 6'h12 ? io_in_1_Re : _GEN_1641; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1649 = _GEN_45 == 6'h12 ? _M0_0_in_waddr_T_2 : _GEN_1644; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1650 = _GEN_45 == 6'h12 ? io_in_2_Im : _GEN_1645; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1651 = _GEN_45 == 6'h12 ? io_in_2_Re : _GEN_1646; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1654 = _GEN_62 == 6'h12 ? _M0_0_in_waddr_T_2 : _GEN_1649; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1655 = _GEN_62 == 6'h12 ? io_in_3_Im : _GEN_1650; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1656 = _GEN_62 == 6'h12 ? io_in_3_Re : _GEN_1651; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1659 = _GEN_79 == 6'h12 ? _M0_0_in_waddr_T_2 : _GEN_1654; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1660 = _GEN_79 == 6'h12 ? io_in_4_Im : _GEN_1655; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1661 = _GEN_79 == 6'h12 ? io_in_4_Re : _GEN_1656; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1664 = _GEN_96 == 6'h12 ? _M0_0_in_waddr_T_2 : _GEN_1659; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1665 = _GEN_96 == 6'h12 ? io_in_5_Im : _GEN_1660; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1666 = _GEN_96 == 6'h12 ? io_in_5_Re : _GEN_1661; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1669 = _GEN_113 == 6'h12 ? _M0_0_in_waddr_T_2 : _GEN_1664; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1670 = _GEN_113 == 6'h12 ? io_in_6_Im : _GEN_1665; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1671 = _GEN_113 == 6'h12 ? io_in_6_Re : _GEN_1666; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1674 = _GEN_130 == 6'h12 ? _M0_0_in_waddr_T_2 : _GEN_1669; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1675 = _GEN_130 == 6'h12 ? io_in_7_Im : _GEN_1670; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1676 = _GEN_130 == 6'h12 ? io_in_7_Re : _GEN_1671; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1679 = _GEN_147 == 6'h12 ? _M0_0_in_waddr_T_26 : _GEN_1674; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1680 = _GEN_147 == 6'h12 ? io_in_8_Im : _GEN_1675; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1681 = _GEN_147 == 6'h12 ? io_in_8_Re : _GEN_1676; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1684 = _GEN_164 == 6'h12 ? _M0_0_in_waddr_T_26 : _GEN_1679; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1685 = _GEN_164 == 6'h12 ? io_in_9_Im : _GEN_1680; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1686 = _GEN_164 == 6'h12 ? io_in_9_Re : _GEN_1681; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1689 = _GEN_181 == 6'h12 ? _M0_0_in_waddr_T_26 : _GEN_1684; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1690 = _GEN_181 == 6'h12 ? io_in_10_Im : _GEN_1685; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1691 = _GEN_181 == 6'h12 ? io_in_10_Re : _GEN_1686; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1694 = _GEN_198 == 6'h12 ? _M0_0_in_waddr_T_26 : _GEN_1689; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1695 = _GEN_198 == 6'h12 ? io_in_11_Im : _GEN_1690; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1696 = _GEN_198 == 6'h12 ? io_in_11_Re : _GEN_1691; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1699 = _GEN_215 == 6'h12 ? _M0_0_in_waddr_T_26 : _GEN_1694; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1700 = _GEN_215 == 6'h12 ? io_in_12_Im : _GEN_1695; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1701 = _GEN_215 == 6'h12 ? io_in_12_Re : _GEN_1696; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1704 = _GEN_232 == 6'h12 ? _M0_0_in_waddr_T_26 : _GEN_1699; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1705 = _GEN_232 == 6'h12 ? io_in_13_Im : _GEN_1700; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1706 = _GEN_232 == 6'h12 ? io_in_13_Re : _GEN_1701; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1708 = _GEN_249 == 6'h12 | (_GEN_232 == 6'h12 | (_GEN_215 == 6'h12 | (_GEN_198 == 6'h12 | (_GEN_181 == 6'h12
     | (_GEN_164 == 6'h12 | (_GEN_147 == 6'h12 | (_GEN_130 == 6'h12 | (_GEN_113 == 6'h12 | (_GEN_96 == 6'h12 | (_GEN_79
     == 6'h12 | (_GEN_62 == 6'h12 | (_GEN_45 == 6'h12 | (_GEN_28 == 6'h12 | _GEN_11 == 6'h12))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1709 = _GEN_249 == 6'h12 ? _M0_0_in_waddr_T_26 : _GEN_1704; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1710 = _GEN_249 == 6'h12 ? io_in_14_Im : _GEN_1705; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1711 = _GEN_249 == 6'h12 ? io_in_14_Re : _GEN_1706; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1713 = _GEN_266 == 6'h12 | _GEN_1708; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1714 = _GEN_266 == 6'h12 ? _M0_0_in_waddr_T_26 : _GEN_1709; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1715 = _GEN_266 == 6'h12 ? io_in_15_Im : _GEN_1710; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1716 = _GEN_266 == 6'h12 ? io_in_15_Re : _GEN_1711; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1719 = _GEN_11 == 6'h13 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1720 = _GEN_11 == 6'h13 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1721 = _GEN_11 == 6'h13 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1724 = _GEN_28 == 6'h13 ? _M0_0_in_waddr_T_2 : _GEN_1719; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1725 = _GEN_28 == 6'h13 ? io_in_1_Im : _GEN_1720; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1726 = _GEN_28 == 6'h13 ? io_in_1_Re : _GEN_1721; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1729 = _GEN_45 == 6'h13 ? _M0_0_in_waddr_T_2 : _GEN_1724; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1730 = _GEN_45 == 6'h13 ? io_in_2_Im : _GEN_1725; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1731 = _GEN_45 == 6'h13 ? io_in_2_Re : _GEN_1726; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1734 = _GEN_62 == 6'h13 ? _M0_0_in_waddr_T_2 : _GEN_1729; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1735 = _GEN_62 == 6'h13 ? io_in_3_Im : _GEN_1730; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1736 = _GEN_62 == 6'h13 ? io_in_3_Re : _GEN_1731; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1739 = _GEN_79 == 6'h13 ? _M0_0_in_waddr_T_2 : _GEN_1734; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1740 = _GEN_79 == 6'h13 ? io_in_4_Im : _GEN_1735; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1741 = _GEN_79 == 6'h13 ? io_in_4_Re : _GEN_1736; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1744 = _GEN_96 == 6'h13 ? _M0_0_in_waddr_T_2 : _GEN_1739; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1745 = _GEN_96 == 6'h13 ? io_in_5_Im : _GEN_1740; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1746 = _GEN_96 == 6'h13 ? io_in_5_Re : _GEN_1741; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1749 = _GEN_113 == 6'h13 ? _M0_0_in_waddr_T_2 : _GEN_1744; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1750 = _GEN_113 == 6'h13 ? io_in_6_Im : _GEN_1745; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1751 = _GEN_113 == 6'h13 ? io_in_6_Re : _GEN_1746; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1754 = _GEN_130 == 6'h13 ? _M0_0_in_waddr_T_2 : _GEN_1749; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1755 = _GEN_130 == 6'h13 ? io_in_7_Im : _GEN_1750; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1756 = _GEN_130 == 6'h13 ? io_in_7_Re : _GEN_1751; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1759 = _GEN_147 == 6'h13 ? _M0_0_in_waddr_T_26 : _GEN_1754; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1760 = _GEN_147 == 6'h13 ? io_in_8_Im : _GEN_1755; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1761 = _GEN_147 == 6'h13 ? io_in_8_Re : _GEN_1756; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1764 = _GEN_164 == 6'h13 ? _M0_0_in_waddr_T_26 : _GEN_1759; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1765 = _GEN_164 == 6'h13 ? io_in_9_Im : _GEN_1760; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1766 = _GEN_164 == 6'h13 ? io_in_9_Re : _GEN_1761; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1769 = _GEN_181 == 6'h13 ? _M0_0_in_waddr_T_26 : _GEN_1764; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1770 = _GEN_181 == 6'h13 ? io_in_10_Im : _GEN_1765; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1771 = _GEN_181 == 6'h13 ? io_in_10_Re : _GEN_1766; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1774 = _GEN_198 == 6'h13 ? _M0_0_in_waddr_T_26 : _GEN_1769; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1775 = _GEN_198 == 6'h13 ? io_in_11_Im : _GEN_1770; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1776 = _GEN_198 == 6'h13 ? io_in_11_Re : _GEN_1771; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1779 = _GEN_215 == 6'h13 ? _M0_0_in_waddr_T_26 : _GEN_1774; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1780 = _GEN_215 == 6'h13 ? io_in_12_Im : _GEN_1775; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1781 = _GEN_215 == 6'h13 ? io_in_12_Re : _GEN_1776; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1784 = _GEN_232 == 6'h13 ? _M0_0_in_waddr_T_26 : _GEN_1779; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1785 = _GEN_232 == 6'h13 ? io_in_13_Im : _GEN_1780; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1786 = _GEN_232 == 6'h13 ? io_in_13_Re : _GEN_1781; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1788 = _GEN_249 == 6'h13 | (_GEN_232 == 6'h13 | (_GEN_215 == 6'h13 | (_GEN_198 == 6'h13 | (_GEN_181 == 6'h13
     | (_GEN_164 == 6'h13 | (_GEN_147 == 6'h13 | (_GEN_130 == 6'h13 | (_GEN_113 == 6'h13 | (_GEN_96 == 6'h13 | (_GEN_79
     == 6'h13 | (_GEN_62 == 6'h13 | (_GEN_45 == 6'h13 | (_GEN_28 == 6'h13 | _GEN_11 == 6'h13))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1789 = _GEN_249 == 6'h13 ? _M0_0_in_waddr_T_26 : _GEN_1784; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1790 = _GEN_249 == 6'h13 ? io_in_14_Im : _GEN_1785; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1791 = _GEN_249 == 6'h13 ? io_in_14_Re : _GEN_1786; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1793 = _GEN_266 == 6'h13 | _GEN_1788; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1794 = _GEN_266 == 6'h13 ? _M0_0_in_waddr_T_26 : _GEN_1789; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1795 = _GEN_266 == 6'h13 ? io_in_15_Im : _GEN_1790; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1796 = _GEN_266 == 6'h13 ? io_in_15_Re : _GEN_1791; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1799 = _GEN_11 == 6'h14 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1800 = _GEN_11 == 6'h14 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1801 = _GEN_11 == 6'h14 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1804 = _GEN_28 == 6'h14 ? _M0_0_in_waddr_T_2 : _GEN_1799; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1805 = _GEN_28 == 6'h14 ? io_in_1_Im : _GEN_1800; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1806 = _GEN_28 == 6'h14 ? io_in_1_Re : _GEN_1801; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1809 = _GEN_45 == 6'h14 ? _M0_0_in_waddr_T_2 : _GEN_1804; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1810 = _GEN_45 == 6'h14 ? io_in_2_Im : _GEN_1805; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1811 = _GEN_45 == 6'h14 ? io_in_2_Re : _GEN_1806; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1814 = _GEN_62 == 6'h14 ? _M0_0_in_waddr_T_2 : _GEN_1809; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1815 = _GEN_62 == 6'h14 ? io_in_3_Im : _GEN_1810; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1816 = _GEN_62 == 6'h14 ? io_in_3_Re : _GEN_1811; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1819 = _GEN_79 == 6'h14 ? _M0_0_in_waddr_T_2 : _GEN_1814; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1820 = _GEN_79 == 6'h14 ? io_in_4_Im : _GEN_1815; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1821 = _GEN_79 == 6'h14 ? io_in_4_Re : _GEN_1816; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1824 = _GEN_96 == 6'h14 ? _M0_0_in_waddr_T_2 : _GEN_1819; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1825 = _GEN_96 == 6'h14 ? io_in_5_Im : _GEN_1820; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1826 = _GEN_96 == 6'h14 ? io_in_5_Re : _GEN_1821; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1829 = _GEN_113 == 6'h14 ? _M0_0_in_waddr_T_2 : _GEN_1824; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1830 = _GEN_113 == 6'h14 ? io_in_6_Im : _GEN_1825; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1831 = _GEN_113 == 6'h14 ? io_in_6_Re : _GEN_1826; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1834 = _GEN_130 == 6'h14 ? _M0_0_in_waddr_T_2 : _GEN_1829; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1835 = _GEN_130 == 6'h14 ? io_in_7_Im : _GEN_1830; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1836 = _GEN_130 == 6'h14 ? io_in_7_Re : _GEN_1831; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1839 = _GEN_147 == 6'h14 ? _M0_0_in_waddr_T_26 : _GEN_1834; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1840 = _GEN_147 == 6'h14 ? io_in_8_Im : _GEN_1835; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1841 = _GEN_147 == 6'h14 ? io_in_8_Re : _GEN_1836; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1844 = _GEN_164 == 6'h14 ? _M0_0_in_waddr_T_26 : _GEN_1839; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1845 = _GEN_164 == 6'h14 ? io_in_9_Im : _GEN_1840; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1846 = _GEN_164 == 6'h14 ? io_in_9_Re : _GEN_1841; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1849 = _GEN_181 == 6'h14 ? _M0_0_in_waddr_T_26 : _GEN_1844; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1850 = _GEN_181 == 6'h14 ? io_in_10_Im : _GEN_1845; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1851 = _GEN_181 == 6'h14 ? io_in_10_Re : _GEN_1846; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1854 = _GEN_198 == 6'h14 ? _M0_0_in_waddr_T_26 : _GEN_1849; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1855 = _GEN_198 == 6'h14 ? io_in_11_Im : _GEN_1850; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1856 = _GEN_198 == 6'h14 ? io_in_11_Re : _GEN_1851; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1859 = _GEN_215 == 6'h14 ? _M0_0_in_waddr_T_26 : _GEN_1854; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1860 = _GEN_215 == 6'h14 ? io_in_12_Im : _GEN_1855; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1861 = _GEN_215 == 6'h14 ? io_in_12_Re : _GEN_1856; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1864 = _GEN_232 == 6'h14 ? _M0_0_in_waddr_T_26 : _GEN_1859; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1865 = _GEN_232 == 6'h14 ? io_in_13_Im : _GEN_1860; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1866 = _GEN_232 == 6'h14 ? io_in_13_Re : _GEN_1861; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1868 = _GEN_249 == 6'h14 | (_GEN_232 == 6'h14 | (_GEN_215 == 6'h14 | (_GEN_198 == 6'h14 | (_GEN_181 == 6'h14
     | (_GEN_164 == 6'h14 | (_GEN_147 == 6'h14 | (_GEN_130 == 6'h14 | (_GEN_113 == 6'h14 | (_GEN_96 == 6'h14 | (_GEN_79
     == 6'h14 | (_GEN_62 == 6'h14 | (_GEN_45 == 6'h14 | (_GEN_28 == 6'h14 | _GEN_11 == 6'h14))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1869 = _GEN_249 == 6'h14 ? _M0_0_in_waddr_T_26 : _GEN_1864; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1870 = _GEN_249 == 6'h14 ? io_in_14_Im : _GEN_1865; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1871 = _GEN_249 == 6'h14 ? io_in_14_Re : _GEN_1866; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1873 = _GEN_266 == 6'h14 | _GEN_1868; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1874 = _GEN_266 == 6'h14 ? _M0_0_in_waddr_T_26 : _GEN_1869; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1875 = _GEN_266 == 6'h14 ? io_in_15_Im : _GEN_1870; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1876 = _GEN_266 == 6'h14 ? io_in_15_Re : _GEN_1871; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1879 = _GEN_11 == 6'h15 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1880 = _GEN_11 == 6'h15 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1881 = _GEN_11 == 6'h15 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1884 = _GEN_28 == 6'h15 ? _M0_0_in_waddr_T_2 : _GEN_1879; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1885 = _GEN_28 == 6'h15 ? io_in_1_Im : _GEN_1880; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1886 = _GEN_28 == 6'h15 ? io_in_1_Re : _GEN_1881; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1889 = _GEN_45 == 6'h15 ? _M0_0_in_waddr_T_2 : _GEN_1884; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1890 = _GEN_45 == 6'h15 ? io_in_2_Im : _GEN_1885; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1891 = _GEN_45 == 6'h15 ? io_in_2_Re : _GEN_1886; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1894 = _GEN_62 == 6'h15 ? _M0_0_in_waddr_T_2 : _GEN_1889; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1895 = _GEN_62 == 6'h15 ? io_in_3_Im : _GEN_1890; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1896 = _GEN_62 == 6'h15 ? io_in_3_Re : _GEN_1891; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1899 = _GEN_79 == 6'h15 ? _M0_0_in_waddr_T_2 : _GEN_1894; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1900 = _GEN_79 == 6'h15 ? io_in_4_Im : _GEN_1895; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1901 = _GEN_79 == 6'h15 ? io_in_4_Re : _GEN_1896; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1904 = _GEN_96 == 6'h15 ? _M0_0_in_waddr_T_2 : _GEN_1899; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1905 = _GEN_96 == 6'h15 ? io_in_5_Im : _GEN_1900; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1906 = _GEN_96 == 6'h15 ? io_in_5_Re : _GEN_1901; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1909 = _GEN_113 == 6'h15 ? _M0_0_in_waddr_T_2 : _GEN_1904; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1910 = _GEN_113 == 6'h15 ? io_in_6_Im : _GEN_1905; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1911 = _GEN_113 == 6'h15 ? io_in_6_Re : _GEN_1906; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1914 = _GEN_130 == 6'h15 ? _M0_0_in_waddr_T_2 : _GEN_1909; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1915 = _GEN_130 == 6'h15 ? io_in_7_Im : _GEN_1910; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1916 = _GEN_130 == 6'h15 ? io_in_7_Re : _GEN_1911; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1919 = _GEN_147 == 6'h15 ? _M0_0_in_waddr_T_26 : _GEN_1914; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1920 = _GEN_147 == 6'h15 ? io_in_8_Im : _GEN_1915; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1921 = _GEN_147 == 6'h15 ? io_in_8_Re : _GEN_1916; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1924 = _GEN_164 == 6'h15 ? _M0_0_in_waddr_T_26 : _GEN_1919; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1925 = _GEN_164 == 6'h15 ? io_in_9_Im : _GEN_1920; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1926 = _GEN_164 == 6'h15 ? io_in_9_Re : _GEN_1921; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1929 = _GEN_181 == 6'h15 ? _M0_0_in_waddr_T_26 : _GEN_1924; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1930 = _GEN_181 == 6'h15 ? io_in_10_Im : _GEN_1925; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1931 = _GEN_181 == 6'h15 ? io_in_10_Re : _GEN_1926; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1934 = _GEN_198 == 6'h15 ? _M0_0_in_waddr_T_26 : _GEN_1929; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1935 = _GEN_198 == 6'h15 ? io_in_11_Im : _GEN_1930; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1936 = _GEN_198 == 6'h15 ? io_in_11_Re : _GEN_1931; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1939 = _GEN_215 == 6'h15 ? _M0_0_in_waddr_T_26 : _GEN_1934; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1940 = _GEN_215 == 6'h15 ? io_in_12_Im : _GEN_1935; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1941 = _GEN_215 == 6'h15 ? io_in_12_Re : _GEN_1936; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1944 = _GEN_232 == 6'h15 ? _M0_0_in_waddr_T_26 : _GEN_1939; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1945 = _GEN_232 == 6'h15 ? io_in_13_Im : _GEN_1940; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1946 = _GEN_232 == 6'h15 ? io_in_13_Re : _GEN_1941; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1948 = _GEN_249 == 6'h15 | (_GEN_232 == 6'h15 | (_GEN_215 == 6'h15 | (_GEN_198 == 6'h15 | (_GEN_181 == 6'h15
     | (_GEN_164 == 6'h15 | (_GEN_147 == 6'h15 | (_GEN_130 == 6'h15 | (_GEN_113 == 6'h15 | (_GEN_96 == 6'h15 | (_GEN_79
     == 6'h15 | (_GEN_62 == 6'h15 | (_GEN_45 == 6'h15 | (_GEN_28 == 6'h15 | _GEN_11 == 6'h15))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1949 = _GEN_249 == 6'h15 ? _M0_0_in_waddr_T_26 : _GEN_1944; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1950 = _GEN_249 == 6'h15 ? io_in_14_Im : _GEN_1945; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1951 = _GEN_249 == 6'h15 ? io_in_14_Re : _GEN_1946; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_1953 = _GEN_266 == 6'h15 | _GEN_1948; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_1954 = _GEN_266 == 6'h15 ? _M0_0_in_waddr_T_26 : _GEN_1949; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1955 = _GEN_266 == 6'h15 ? io_in_15_Im : _GEN_1950; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1956 = _GEN_266 == 6'h15 ? io_in_15_Re : _GEN_1951; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1959 = _GEN_11 == 6'h16 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_1960 = _GEN_11 == 6'h16 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_1961 = _GEN_11 == 6'h16 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_1964 = _GEN_28 == 6'h16 ? _M0_0_in_waddr_T_2 : _GEN_1959; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1965 = _GEN_28 == 6'h16 ? io_in_1_Im : _GEN_1960; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1966 = _GEN_28 == 6'h16 ? io_in_1_Re : _GEN_1961; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1969 = _GEN_45 == 6'h16 ? _M0_0_in_waddr_T_2 : _GEN_1964; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1970 = _GEN_45 == 6'h16 ? io_in_2_Im : _GEN_1965; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1971 = _GEN_45 == 6'h16 ? io_in_2_Re : _GEN_1966; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1974 = _GEN_62 == 6'h16 ? _M0_0_in_waddr_T_2 : _GEN_1969; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1975 = _GEN_62 == 6'h16 ? io_in_3_Im : _GEN_1970; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1976 = _GEN_62 == 6'h16 ? io_in_3_Re : _GEN_1971; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1979 = _GEN_79 == 6'h16 ? _M0_0_in_waddr_T_2 : _GEN_1974; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1980 = _GEN_79 == 6'h16 ? io_in_4_Im : _GEN_1975; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1981 = _GEN_79 == 6'h16 ? io_in_4_Re : _GEN_1976; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1984 = _GEN_96 == 6'h16 ? _M0_0_in_waddr_T_2 : _GEN_1979; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1985 = _GEN_96 == 6'h16 ? io_in_5_Im : _GEN_1980; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1986 = _GEN_96 == 6'h16 ? io_in_5_Re : _GEN_1981; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1989 = _GEN_113 == 6'h16 ? _M0_0_in_waddr_T_2 : _GEN_1984; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1990 = _GEN_113 == 6'h16 ? io_in_6_Im : _GEN_1985; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1991 = _GEN_113 == 6'h16 ? io_in_6_Re : _GEN_1986; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1994 = _GEN_130 == 6'h16 ? _M0_0_in_waddr_T_2 : _GEN_1989; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_1995 = _GEN_130 == 6'h16 ? io_in_7_Im : _GEN_1990; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_1996 = _GEN_130 == 6'h16 ? io_in_7_Re : _GEN_1991; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_1999 = _GEN_147 == 6'h16 ? _M0_0_in_waddr_T_26 : _GEN_1994; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2000 = _GEN_147 == 6'h16 ? io_in_8_Im : _GEN_1995; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2001 = _GEN_147 == 6'h16 ? io_in_8_Re : _GEN_1996; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2004 = _GEN_164 == 6'h16 ? _M0_0_in_waddr_T_26 : _GEN_1999; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2005 = _GEN_164 == 6'h16 ? io_in_9_Im : _GEN_2000; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2006 = _GEN_164 == 6'h16 ? io_in_9_Re : _GEN_2001; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2009 = _GEN_181 == 6'h16 ? _M0_0_in_waddr_T_26 : _GEN_2004; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2010 = _GEN_181 == 6'h16 ? io_in_10_Im : _GEN_2005; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2011 = _GEN_181 == 6'h16 ? io_in_10_Re : _GEN_2006; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2014 = _GEN_198 == 6'h16 ? _M0_0_in_waddr_T_26 : _GEN_2009; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2015 = _GEN_198 == 6'h16 ? io_in_11_Im : _GEN_2010; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2016 = _GEN_198 == 6'h16 ? io_in_11_Re : _GEN_2011; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2019 = _GEN_215 == 6'h16 ? _M0_0_in_waddr_T_26 : _GEN_2014; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2020 = _GEN_215 == 6'h16 ? io_in_12_Im : _GEN_2015; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2021 = _GEN_215 == 6'h16 ? io_in_12_Re : _GEN_2016; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2024 = _GEN_232 == 6'h16 ? _M0_0_in_waddr_T_26 : _GEN_2019; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2025 = _GEN_232 == 6'h16 ? io_in_13_Im : _GEN_2020; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2026 = _GEN_232 == 6'h16 ? io_in_13_Re : _GEN_2021; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_2028 = _GEN_249 == 6'h16 | (_GEN_232 == 6'h16 | (_GEN_215 == 6'h16 | (_GEN_198 == 6'h16 | (_GEN_181 == 6'h16
     | (_GEN_164 == 6'h16 | (_GEN_147 == 6'h16 | (_GEN_130 == 6'h16 | (_GEN_113 == 6'h16 | (_GEN_96 == 6'h16 | (_GEN_79
     == 6'h16 | (_GEN_62 == 6'h16 | (_GEN_45 == 6'h16 | (_GEN_28 == 6'h16 | _GEN_11 == 6'h16))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_2029 = _GEN_249 == 6'h16 ? _M0_0_in_waddr_T_26 : _GEN_2024; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2030 = _GEN_249 == 6'h16 ? io_in_14_Im : _GEN_2025; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2031 = _GEN_249 == 6'h16 ? io_in_14_Re : _GEN_2026; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_2033 = _GEN_266 == 6'h16 | _GEN_2028; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_2034 = _GEN_266 == 6'h16 ? _M0_0_in_waddr_T_26 : _GEN_2029; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2035 = _GEN_266 == 6'h16 ? io_in_15_Im : _GEN_2030; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2036 = _GEN_266 == 6'h16 ? io_in_15_Re : _GEN_2031; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2039 = _GEN_11 == 6'h17 ? _M0_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2791:26 2797:44 2799:30]
  wire [31:0] _GEN_2040 = _GEN_11 == 6'h17 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [31:0] _GEN_2041 = _GEN_11 == 6'h17 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2792:25 2797:44 2800:29]
  wire [3:0] _GEN_2044 = _GEN_28 == 6'h17 ? _M0_0_in_waddr_T_2 : _GEN_2039; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2045 = _GEN_28 == 6'h17 ? io_in_1_Im : _GEN_2040; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2046 = _GEN_28 == 6'h17 ? io_in_1_Re : _GEN_2041; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2049 = _GEN_45 == 6'h17 ? _M0_0_in_waddr_T_2 : _GEN_2044; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2050 = _GEN_45 == 6'h17 ? io_in_2_Im : _GEN_2045; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2051 = _GEN_45 == 6'h17 ? io_in_2_Re : _GEN_2046; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2054 = _GEN_62 == 6'h17 ? _M0_0_in_waddr_T_2 : _GEN_2049; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2055 = _GEN_62 == 6'h17 ? io_in_3_Im : _GEN_2050; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2056 = _GEN_62 == 6'h17 ? io_in_3_Re : _GEN_2051; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2059 = _GEN_79 == 6'h17 ? _M0_0_in_waddr_T_2 : _GEN_2054; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2060 = _GEN_79 == 6'h17 ? io_in_4_Im : _GEN_2055; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2061 = _GEN_79 == 6'h17 ? io_in_4_Re : _GEN_2056; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2064 = _GEN_96 == 6'h17 ? _M0_0_in_waddr_T_2 : _GEN_2059; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2065 = _GEN_96 == 6'h17 ? io_in_5_Im : _GEN_2060; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2066 = _GEN_96 == 6'h17 ? io_in_5_Re : _GEN_2061; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2069 = _GEN_113 == 6'h17 ? _M0_0_in_waddr_T_2 : _GEN_2064; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2070 = _GEN_113 == 6'h17 ? io_in_6_Im : _GEN_2065; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2071 = _GEN_113 == 6'h17 ? io_in_6_Re : _GEN_2066; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2074 = _GEN_130 == 6'h17 ? _M0_0_in_waddr_T_2 : _GEN_2069; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2075 = _GEN_130 == 6'h17 ? io_in_7_Im : _GEN_2070; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2076 = _GEN_130 == 6'h17 ? io_in_7_Re : _GEN_2071; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2079 = _GEN_147 == 6'h17 ? _M0_0_in_waddr_T_26 : _GEN_2074; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2080 = _GEN_147 == 6'h17 ? io_in_8_Im : _GEN_2075; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2081 = _GEN_147 == 6'h17 ? io_in_8_Re : _GEN_2076; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2084 = _GEN_164 == 6'h17 ? _M0_0_in_waddr_T_26 : _GEN_2079; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2085 = _GEN_164 == 6'h17 ? io_in_9_Im : _GEN_2080; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2086 = _GEN_164 == 6'h17 ? io_in_9_Re : _GEN_2081; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2089 = _GEN_181 == 6'h17 ? _M0_0_in_waddr_T_26 : _GEN_2084; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2090 = _GEN_181 == 6'h17 ? io_in_10_Im : _GEN_2085; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2091 = _GEN_181 == 6'h17 ? io_in_10_Re : _GEN_2086; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2094 = _GEN_198 == 6'h17 ? _M0_0_in_waddr_T_26 : _GEN_2089; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2095 = _GEN_198 == 6'h17 ? io_in_11_Im : _GEN_2090; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2096 = _GEN_198 == 6'h17 ? io_in_11_Re : _GEN_2091; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2099 = _GEN_215 == 6'h17 ? _M0_0_in_waddr_T_26 : _GEN_2094; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2100 = _GEN_215 == 6'h17 ? io_in_12_Im : _GEN_2095; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2101 = _GEN_215 == 6'h17 ? io_in_12_Re : _GEN_2096; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2104 = _GEN_232 == 6'h17 ? _M0_0_in_waddr_T_26 : _GEN_2099; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2105 = _GEN_232 == 6'h17 ? io_in_13_Im : _GEN_2100; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2106 = _GEN_232 == 6'h17 ? io_in_13_Re : _GEN_2101; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_2108 = _GEN_249 == 6'h17 | (_GEN_232 == 6'h17 | (_GEN_215 == 6'h17 | (_GEN_198 == 6'h17 | (_GEN_181 == 6'h17
     | (_GEN_164 == 6'h17 | (_GEN_147 == 6'h17 | (_GEN_130 == 6'h17 | (_GEN_113 == 6'h17 | (_GEN_96 == 6'h17 | (_GEN_79
     == 6'h17 | (_GEN_62 == 6'h17 | (_GEN_45 == 6'h17 | (_GEN_28 == 6'h17 | _GEN_11 == 6'h17))))))))))))); // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_2109 = _GEN_249 == 6'h17 ? _M0_0_in_waddr_T_26 : _GEN_2104; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2110 = _GEN_249 == 6'h17 ? io_in_14_Im : _GEN_2105; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2111 = _GEN_249 == 6'h17 ? io_in_14_Re : _GEN_2106; // @[FFTDesigns.scala 2797:44 2800:29]
  wire  _GEN_2113 = _GEN_266 == 6'h17 | _GEN_2108; // @[FFTDesigns.scala 2797:44 2798:24]
  wire [3:0] _GEN_2114 = _GEN_266 == 6'h17 ? _M0_0_in_waddr_T_26 : _GEN_2109; // @[FFTDesigns.scala 2797:44 2799:30]
  wire [31:0] _GEN_2115 = _GEN_266 == 6'h17 ? io_in_15_Im : _GEN_2110; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [31:0] _GEN_2116 = _GEN_266 == 6'h17 ? io_in_15_Re : _GEN_2111; // @[FFTDesigns.scala 2797:44 2800:29]
  wire [3:0] _GEN_2122 = M0_0_re ? _M0_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2123 = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2781:26 2816:26]
  wire [3:0] _GEN_2124 = M0_0_re ? _M1_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2132 = M0_0_re ? _M0_1_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2134 = M0_0_re ? _M1_1_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2142 = M0_0_re ? _M0_2_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2144 = M0_0_re ? _M1_2_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2152 = M0_0_re ? _M0_3_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2154 = M0_0_re ? _M1_3_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2162 = M0_0_re ? _M0_4_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2164 = M0_0_re ? _M1_4_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2172 = M0_0_re ? _M0_5_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2174 = M0_0_re ? _M1_5_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2182 = M0_0_re ? _M0_6_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2184 = M0_0_re ? _M1_6_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2192 = M0_0_re ? _M0_7_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2194 = M0_0_re ? _M1_7_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2202 = M0_0_re ? _M0_8_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2204 = M0_0_re ? _M1_8_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2212 = M0_0_re ? _M0_9_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2214 = M0_0_re ? _M1_9_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2222 = M0_0_re ? _M0_10_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2224 = M0_0_re ? _M1_10_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2232 = M0_0_re ? _M0_11_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2234 = M0_0_re ? _M1_11_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2242 = M0_0_re ? _M0_12_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2244 = M0_0_re ? _M1_12_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2252 = M0_0_re ? _M0_13_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2254 = M0_0_re ? _M1_13_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2262 = M0_0_re ? _M0_14_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2264 = M0_0_re ? _M1_14_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2272 = M0_0_re ? _M0_15_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2274 = M0_0_re ? _M1_15_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2282 = M0_0_re ? _M0_16_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2284 = M0_0_re ? _M1_16_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2292 = M0_0_re ? _M0_17_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2294 = M0_0_re ? _M1_17_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2302 = M0_0_re ? _M0_18_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2304 = M0_0_re ? _M1_18_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2312 = M0_0_re ? _M0_19_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2314 = M0_0_re ? _M1_19_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2322 = M0_0_re ? _M0_20_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2324 = M0_0_re ? _M1_20_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2332 = M0_0_re ? _M0_21_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2334 = M0_0_re ? _M1_21_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2342 = M0_0_re ? _M0_22_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2344 = M0_0_re ? _M1_22_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2352 = M0_0_re ? _M0_23_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2757:33 2778:26 2813:26]
  wire [3:0] _GEN_2354 = M0_0_re ? _M1_23_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2757:33 2782:26 2817:26]
  wire [3:0] _GEN_2363 = M0_0_re ? _GEN_274 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2368 = M0_0_re ? _GEN_354 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2373 = M0_0_re ? _GEN_434 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2378 = M0_0_re ? _GEN_514 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2383 = M0_0_re ? _GEN_594 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2388 = M0_0_re ? _GEN_674 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2393 = M0_0_re ? _GEN_754 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2398 = M0_0_re ? _GEN_834 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2403 = M0_0_re ? _GEN_914 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2408 = M0_0_re ? _GEN_994 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2413 = M0_0_re ? _GEN_1074 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2418 = M0_0_re ? _GEN_1154 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2423 = M0_0_re ? _GEN_1234 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2428 = M0_0_re ? _GEN_1314 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2433 = M0_0_re ? _GEN_1394 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2438 = M0_0_re ? _GEN_1474 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2443 = M0_0_re ? _GEN_1554 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2448 = M0_0_re ? _GEN_1634 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2453 = M0_0_re ? _GEN_1714 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2458 = M0_0_re ? _GEN_1794 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2463 = M0_0_re ? _GEN_1874 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2468 = M0_0_re ? _GEN_1954 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2473 = M0_0_re ? _GEN_2034 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  wire [3:0] _GEN_2478 = M0_0_re ? _GEN_2114 : 4'h0; // @[FFTDesigns.scala 2757:33 2814:26]
  RAM_Block_224 RAM_Block ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_1 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_2 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_3 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_4 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_5 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_6 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_7 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_8 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_9 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_10 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_11 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_12 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_13 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_14 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_15 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_16 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_16_clock),
    .io_in_raddr(RAM_Block_16_io_in_raddr),
    .io_in_waddr(RAM_Block_16_io_in_waddr),
    .io_in_data_Re(RAM_Block_16_io_in_data_Re),
    .io_in_data_Im(RAM_Block_16_io_in_data_Im),
    .io_re(RAM_Block_16_io_re),
    .io_wr(RAM_Block_16_io_wr),
    .io_en(RAM_Block_16_io_en),
    .io_out_data_Re(RAM_Block_16_io_out_data_Re),
    .io_out_data_Im(RAM_Block_16_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_17 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_17_clock),
    .io_in_raddr(RAM_Block_17_io_in_raddr),
    .io_in_waddr(RAM_Block_17_io_in_waddr),
    .io_in_data_Re(RAM_Block_17_io_in_data_Re),
    .io_in_data_Im(RAM_Block_17_io_in_data_Im),
    .io_re(RAM_Block_17_io_re),
    .io_wr(RAM_Block_17_io_wr),
    .io_en(RAM_Block_17_io_en),
    .io_out_data_Re(RAM_Block_17_io_out_data_Re),
    .io_out_data_Im(RAM_Block_17_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_18 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_18_clock),
    .io_in_raddr(RAM_Block_18_io_in_raddr),
    .io_in_waddr(RAM_Block_18_io_in_waddr),
    .io_in_data_Re(RAM_Block_18_io_in_data_Re),
    .io_in_data_Im(RAM_Block_18_io_in_data_Im),
    .io_re(RAM_Block_18_io_re),
    .io_wr(RAM_Block_18_io_wr),
    .io_en(RAM_Block_18_io_en),
    .io_out_data_Re(RAM_Block_18_io_out_data_Re),
    .io_out_data_Im(RAM_Block_18_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_19 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_19_clock),
    .io_in_raddr(RAM_Block_19_io_in_raddr),
    .io_in_waddr(RAM_Block_19_io_in_waddr),
    .io_in_data_Re(RAM_Block_19_io_in_data_Re),
    .io_in_data_Im(RAM_Block_19_io_in_data_Im),
    .io_re(RAM_Block_19_io_re),
    .io_wr(RAM_Block_19_io_wr),
    .io_en(RAM_Block_19_io_en),
    .io_out_data_Re(RAM_Block_19_io_out_data_Re),
    .io_out_data_Im(RAM_Block_19_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_20 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_20_clock),
    .io_in_raddr(RAM_Block_20_io_in_raddr),
    .io_in_waddr(RAM_Block_20_io_in_waddr),
    .io_in_data_Re(RAM_Block_20_io_in_data_Re),
    .io_in_data_Im(RAM_Block_20_io_in_data_Im),
    .io_re(RAM_Block_20_io_re),
    .io_wr(RAM_Block_20_io_wr),
    .io_en(RAM_Block_20_io_en),
    .io_out_data_Re(RAM_Block_20_io_out_data_Re),
    .io_out_data_Im(RAM_Block_20_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_21 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_21_clock),
    .io_in_raddr(RAM_Block_21_io_in_raddr),
    .io_in_waddr(RAM_Block_21_io_in_waddr),
    .io_in_data_Re(RAM_Block_21_io_in_data_Re),
    .io_in_data_Im(RAM_Block_21_io_in_data_Im),
    .io_re(RAM_Block_21_io_re),
    .io_wr(RAM_Block_21_io_wr),
    .io_en(RAM_Block_21_io_en),
    .io_out_data_Re(RAM_Block_21_io_out_data_Re),
    .io_out_data_Im(RAM_Block_21_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_22 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_22_clock),
    .io_in_raddr(RAM_Block_22_io_in_raddr),
    .io_in_waddr(RAM_Block_22_io_in_waddr),
    .io_in_data_Re(RAM_Block_22_io_in_data_Re),
    .io_in_data_Im(RAM_Block_22_io_in_data_Im),
    .io_re(RAM_Block_22_io_re),
    .io_wr(RAM_Block_22_io_wr),
    .io_en(RAM_Block_22_io_en),
    .io_out_data_Re(RAM_Block_22_io_out_data_Re),
    .io_out_data_Im(RAM_Block_22_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_23 ( // @[FFTDesigns.scala 2713:26]
    .clock(RAM_Block_23_clock),
    .io_in_raddr(RAM_Block_23_io_in_raddr),
    .io_in_waddr(RAM_Block_23_io_in_waddr),
    .io_in_data_Re(RAM_Block_23_io_in_data_Re),
    .io_in_data_Im(RAM_Block_23_io_in_data_Im),
    .io_re(RAM_Block_23_io_re),
    .io_wr(RAM_Block_23_io_wr),
    .io_en(RAM_Block_23_io_en),
    .io_out_data_Re(RAM_Block_23_io_out_data_Re),
    .io_out_data_Im(RAM_Block_23_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_24 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_24_clock),
    .io_in_raddr(RAM_Block_24_io_in_raddr),
    .io_in_waddr(RAM_Block_24_io_in_waddr),
    .io_in_data_Re(RAM_Block_24_io_in_data_Re),
    .io_in_data_Im(RAM_Block_24_io_in_data_Im),
    .io_re(RAM_Block_24_io_re),
    .io_wr(RAM_Block_24_io_wr),
    .io_en(RAM_Block_24_io_en),
    .io_out_data_Re(RAM_Block_24_io_out_data_Re),
    .io_out_data_Im(RAM_Block_24_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_25 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_25_clock),
    .io_in_raddr(RAM_Block_25_io_in_raddr),
    .io_in_waddr(RAM_Block_25_io_in_waddr),
    .io_in_data_Re(RAM_Block_25_io_in_data_Re),
    .io_in_data_Im(RAM_Block_25_io_in_data_Im),
    .io_re(RAM_Block_25_io_re),
    .io_wr(RAM_Block_25_io_wr),
    .io_en(RAM_Block_25_io_en),
    .io_out_data_Re(RAM_Block_25_io_out_data_Re),
    .io_out_data_Im(RAM_Block_25_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_26 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_26_clock),
    .io_in_raddr(RAM_Block_26_io_in_raddr),
    .io_in_waddr(RAM_Block_26_io_in_waddr),
    .io_in_data_Re(RAM_Block_26_io_in_data_Re),
    .io_in_data_Im(RAM_Block_26_io_in_data_Im),
    .io_re(RAM_Block_26_io_re),
    .io_wr(RAM_Block_26_io_wr),
    .io_en(RAM_Block_26_io_en),
    .io_out_data_Re(RAM_Block_26_io_out_data_Re),
    .io_out_data_Im(RAM_Block_26_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_27 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_27_clock),
    .io_in_raddr(RAM_Block_27_io_in_raddr),
    .io_in_waddr(RAM_Block_27_io_in_waddr),
    .io_in_data_Re(RAM_Block_27_io_in_data_Re),
    .io_in_data_Im(RAM_Block_27_io_in_data_Im),
    .io_re(RAM_Block_27_io_re),
    .io_wr(RAM_Block_27_io_wr),
    .io_en(RAM_Block_27_io_en),
    .io_out_data_Re(RAM_Block_27_io_out_data_Re),
    .io_out_data_Im(RAM_Block_27_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_28 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_28_clock),
    .io_in_raddr(RAM_Block_28_io_in_raddr),
    .io_in_waddr(RAM_Block_28_io_in_waddr),
    .io_in_data_Re(RAM_Block_28_io_in_data_Re),
    .io_in_data_Im(RAM_Block_28_io_in_data_Im),
    .io_re(RAM_Block_28_io_re),
    .io_wr(RAM_Block_28_io_wr),
    .io_en(RAM_Block_28_io_en),
    .io_out_data_Re(RAM_Block_28_io_out_data_Re),
    .io_out_data_Im(RAM_Block_28_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_29 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_29_clock),
    .io_in_raddr(RAM_Block_29_io_in_raddr),
    .io_in_waddr(RAM_Block_29_io_in_waddr),
    .io_in_data_Re(RAM_Block_29_io_in_data_Re),
    .io_in_data_Im(RAM_Block_29_io_in_data_Im),
    .io_re(RAM_Block_29_io_re),
    .io_wr(RAM_Block_29_io_wr),
    .io_en(RAM_Block_29_io_en),
    .io_out_data_Re(RAM_Block_29_io_out_data_Re),
    .io_out_data_Im(RAM_Block_29_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_30 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_30_clock),
    .io_in_raddr(RAM_Block_30_io_in_raddr),
    .io_in_waddr(RAM_Block_30_io_in_waddr),
    .io_in_data_Re(RAM_Block_30_io_in_data_Re),
    .io_in_data_Im(RAM_Block_30_io_in_data_Im),
    .io_re(RAM_Block_30_io_re),
    .io_wr(RAM_Block_30_io_wr),
    .io_en(RAM_Block_30_io_en),
    .io_out_data_Re(RAM_Block_30_io_out_data_Re),
    .io_out_data_Im(RAM_Block_30_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_31 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_31_clock),
    .io_in_raddr(RAM_Block_31_io_in_raddr),
    .io_in_waddr(RAM_Block_31_io_in_waddr),
    .io_in_data_Re(RAM_Block_31_io_in_data_Re),
    .io_in_data_Im(RAM_Block_31_io_in_data_Im),
    .io_re(RAM_Block_31_io_re),
    .io_wr(RAM_Block_31_io_wr),
    .io_en(RAM_Block_31_io_en),
    .io_out_data_Re(RAM_Block_31_io_out_data_Re),
    .io_out_data_Im(RAM_Block_31_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_32 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_32_clock),
    .io_in_raddr(RAM_Block_32_io_in_raddr),
    .io_in_waddr(RAM_Block_32_io_in_waddr),
    .io_in_data_Re(RAM_Block_32_io_in_data_Re),
    .io_in_data_Im(RAM_Block_32_io_in_data_Im),
    .io_re(RAM_Block_32_io_re),
    .io_wr(RAM_Block_32_io_wr),
    .io_en(RAM_Block_32_io_en),
    .io_out_data_Re(RAM_Block_32_io_out_data_Re),
    .io_out_data_Im(RAM_Block_32_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_33 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_33_clock),
    .io_in_raddr(RAM_Block_33_io_in_raddr),
    .io_in_waddr(RAM_Block_33_io_in_waddr),
    .io_in_data_Re(RAM_Block_33_io_in_data_Re),
    .io_in_data_Im(RAM_Block_33_io_in_data_Im),
    .io_re(RAM_Block_33_io_re),
    .io_wr(RAM_Block_33_io_wr),
    .io_en(RAM_Block_33_io_en),
    .io_out_data_Re(RAM_Block_33_io_out_data_Re),
    .io_out_data_Im(RAM_Block_33_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_34 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_34_clock),
    .io_in_raddr(RAM_Block_34_io_in_raddr),
    .io_in_waddr(RAM_Block_34_io_in_waddr),
    .io_in_data_Re(RAM_Block_34_io_in_data_Re),
    .io_in_data_Im(RAM_Block_34_io_in_data_Im),
    .io_re(RAM_Block_34_io_re),
    .io_wr(RAM_Block_34_io_wr),
    .io_en(RAM_Block_34_io_en),
    .io_out_data_Re(RAM_Block_34_io_out_data_Re),
    .io_out_data_Im(RAM_Block_34_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_35 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_35_clock),
    .io_in_raddr(RAM_Block_35_io_in_raddr),
    .io_in_waddr(RAM_Block_35_io_in_waddr),
    .io_in_data_Re(RAM_Block_35_io_in_data_Re),
    .io_in_data_Im(RAM_Block_35_io_in_data_Im),
    .io_re(RAM_Block_35_io_re),
    .io_wr(RAM_Block_35_io_wr),
    .io_en(RAM_Block_35_io_en),
    .io_out_data_Re(RAM_Block_35_io_out_data_Re),
    .io_out_data_Im(RAM_Block_35_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_36 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_36_clock),
    .io_in_raddr(RAM_Block_36_io_in_raddr),
    .io_in_waddr(RAM_Block_36_io_in_waddr),
    .io_in_data_Re(RAM_Block_36_io_in_data_Re),
    .io_in_data_Im(RAM_Block_36_io_in_data_Im),
    .io_re(RAM_Block_36_io_re),
    .io_wr(RAM_Block_36_io_wr),
    .io_en(RAM_Block_36_io_en),
    .io_out_data_Re(RAM_Block_36_io_out_data_Re),
    .io_out_data_Im(RAM_Block_36_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_37 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_37_clock),
    .io_in_raddr(RAM_Block_37_io_in_raddr),
    .io_in_waddr(RAM_Block_37_io_in_waddr),
    .io_in_data_Re(RAM_Block_37_io_in_data_Re),
    .io_in_data_Im(RAM_Block_37_io_in_data_Im),
    .io_re(RAM_Block_37_io_re),
    .io_wr(RAM_Block_37_io_wr),
    .io_en(RAM_Block_37_io_en),
    .io_out_data_Re(RAM_Block_37_io_out_data_Re),
    .io_out_data_Im(RAM_Block_37_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_38 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_38_clock),
    .io_in_raddr(RAM_Block_38_io_in_raddr),
    .io_in_waddr(RAM_Block_38_io_in_waddr),
    .io_in_data_Re(RAM_Block_38_io_in_data_Re),
    .io_in_data_Im(RAM_Block_38_io_in_data_Im),
    .io_re(RAM_Block_38_io_re),
    .io_wr(RAM_Block_38_io_wr),
    .io_en(RAM_Block_38_io_en),
    .io_out_data_Re(RAM_Block_38_io_out_data_Re),
    .io_out_data_Im(RAM_Block_38_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_39 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_39_clock),
    .io_in_raddr(RAM_Block_39_io_in_raddr),
    .io_in_waddr(RAM_Block_39_io_in_waddr),
    .io_in_data_Re(RAM_Block_39_io_in_data_Re),
    .io_in_data_Im(RAM_Block_39_io_in_data_Im),
    .io_re(RAM_Block_39_io_re),
    .io_wr(RAM_Block_39_io_wr),
    .io_en(RAM_Block_39_io_en),
    .io_out_data_Re(RAM_Block_39_io_out_data_Re),
    .io_out_data_Im(RAM_Block_39_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_40 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_40_clock),
    .io_in_raddr(RAM_Block_40_io_in_raddr),
    .io_in_waddr(RAM_Block_40_io_in_waddr),
    .io_in_data_Re(RAM_Block_40_io_in_data_Re),
    .io_in_data_Im(RAM_Block_40_io_in_data_Im),
    .io_re(RAM_Block_40_io_re),
    .io_wr(RAM_Block_40_io_wr),
    .io_en(RAM_Block_40_io_en),
    .io_out_data_Re(RAM_Block_40_io_out_data_Re),
    .io_out_data_Im(RAM_Block_40_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_41 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_41_clock),
    .io_in_raddr(RAM_Block_41_io_in_raddr),
    .io_in_waddr(RAM_Block_41_io_in_waddr),
    .io_in_data_Re(RAM_Block_41_io_in_data_Re),
    .io_in_data_Im(RAM_Block_41_io_in_data_Im),
    .io_re(RAM_Block_41_io_re),
    .io_wr(RAM_Block_41_io_wr),
    .io_en(RAM_Block_41_io_en),
    .io_out_data_Re(RAM_Block_41_io_out_data_Re),
    .io_out_data_Im(RAM_Block_41_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_42 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_42_clock),
    .io_in_raddr(RAM_Block_42_io_in_raddr),
    .io_in_waddr(RAM_Block_42_io_in_waddr),
    .io_in_data_Re(RAM_Block_42_io_in_data_Re),
    .io_in_data_Im(RAM_Block_42_io_in_data_Im),
    .io_re(RAM_Block_42_io_re),
    .io_wr(RAM_Block_42_io_wr),
    .io_en(RAM_Block_42_io_en),
    .io_out_data_Re(RAM_Block_42_io_out_data_Re),
    .io_out_data_Im(RAM_Block_42_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_43 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_43_clock),
    .io_in_raddr(RAM_Block_43_io_in_raddr),
    .io_in_waddr(RAM_Block_43_io_in_waddr),
    .io_in_data_Re(RAM_Block_43_io_in_data_Re),
    .io_in_data_Im(RAM_Block_43_io_in_data_Im),
    .io_re(RAM_Block_43_io_re),
    .io_wr(RAM_Block_43_io_wr),
    .io_en(RAM_Block_43_io_en),
    .io_out_data_Re(RAM_Block_43_io_out_data_Re),
    .io_out_data_Im(RAM_Block_43_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_44 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_44_clock),
    .io_in_raddr(RAM_Block_44_io_in_raddr),
    .io_in_waddr(RAM_Block_44_io_in_waddr),
    .io_in_data_Re(RAM_Block_44_io_in_data_Re),
    .io_in_data_Im(RAM_Block_44_io_in_data_Im),
    .io_re(RAM_Block_44_io_re),
    .io_wr(RAM_Block_44_io_wr),
    .io_en(RAM_Block_44_io_en),
    .io_out_data_Re(RAM_Block_44_io_out_data_Re),
    .io_out_data_Im(RAM_Block_44_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_45 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_45_clock),
    .io_in_raddr(RAM_Block_45_io_in_raddr),
    .io_in_waddr(RAM_Block_45_io_in_waddr),
    .io_in_data_Re(RAM_Block_45_io_in_data_Re),
    .io_in_data_Im(RAM_Block_45_io_in_data_Im),
    .io_re(RAM_Block_45_io_re),
    .io_wr(RAM_Block_45_io_wr),
    .io_en(RAM_Block_45_io_en),
    .io_out_data_Re(RAM_Block_45_io_out_data_Re),
    .io_out_data_Im(RAM_Block_45_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_46 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_46_clock),
    .io_in_raddr(RAM_Block_46_io_in_raddr),
    .io_in_waddr(RAM_Block_46_io_in_waddr),
    .io_in_data_Re(RAM_Block_46_io_in_data_Re),
    .io_in_data_Im(RAM_Block_46_io_in_data_Im),
    .io_re(RAM_Block_46_io_re),
    .io_wr(RAM_Block_46_io_wr),
    .io_en(RAM_Block_46_io_en),
    .io_out_data_Re(RAM_Block_46_io_out_data_Re),
    .io_out_data_Im(RAM_Block_46_io_out_data_Im)
  );
  RAM_Block_224 RAM_Block_47 ( // @[FFTDesigns.scala 2717:26]
    .clock(RAM_Block_47_clock),
    .io_in_raddr(RAM_Block_47_io_in_raddr),
    .io_in_waddr(RAM_Block_47_io_in_waddr),
    .io_in_data_Re(RAM_Block_47_io_in_data_Re),
    .io_in_data_Im(RAM_Block_47_io_in_data_Im),
    .io_re(RAM_Block_47_io_re),
    .io_wr(RAM_Block_47_io_wr),
    .io_en(RAM_Block_47_io_en),
    .io_out_data_Re(RAM_Block_47_io_out_data_Re),
    .io_out_data_Im(RAM_Block_47_io_out_data_Im)
  );
  PermutationModuleStreamed_7 PermutationModuleStreamed ( // @[FFTDesigns.scala 2750:28]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_8_Re(PermutationModuleStreamed_io_in_8_Re),
    .io_in_8_Im(PermutationModuleStreamed_io_in_8_Im),
    .io_in_9_Re(PermutationModuleStreamed_io_in_9_Re),
    .io_in_9_Im(PermutationModuleStreamed_io_in_9_Im),
    .io_in_10_Re(PermutationModuleStreamed_io_in_10_Re),
    .io_in_10_Im(PermutationModuleStreamed_io_in_10_Im),
    .io_in_11_Re(PermutationModuleStreamed_io_in_11_Re),
    .io_in_11_Im(PermutationModuleStreamed_io_in_11_Im),
    .io_in_12_Re(PermutationModuleStreamed_io_in_12_Re),
    .io_in_12_Im(PermutationModuleStreamed_io_in_12_Im),
    .io_in_13_Re(PermutationModuleStreamed_io_in_13_Re),
    .io_in_13_Im(PermutationModuleStreamed_io_in_13_Im),
    .io_in_14_Re(PermutationModuleStreamed_io_in_14_Re),
    .io_in_14_Im(PermutationModuleStreamed_io_in_14_Im),
    .io_in_15_Re(PermutationModuleStreamed_io_in_15_Re),
    .io_in_15_Im(PermutationModuleStreamed_io_in_15_Im),
    .io_in_16_Re(PermutationModuleStreamed_io_in_16_Re),
    .io_in_16_Im(PermutationModuleStreamed_io_in_16_Im),
    .io_in_17_Re(PermutationModuleStreamed_io_in_17_Re),
    .io_in_17_Im(PermutationModuleStreamed_io_in_17_Im),
    .io_in_18_Re(PermutationModuleStreamed_io_in_18_Re),
    .io_in_18_Im(PermutationModuleStreamed_io_in_18_Im),
    .io_in_19_Re(PermutationModuleStreamed_io_in_19_Re),
    .io_in_19_Im(PermutationModuleStreamed_io_in_19_Im),
    .io_in_20_Re(PermutationModuleStreamed_io_in_20_Re),
    .io_in_20_Im(PermutationModuleStreamed_io_in_20_Im),
    .io_in_21_Re(PermutationModuleStreamed_io_in_21_Re),
    .io_in_21_Im(PermutationModuleStreamed_io_in_21_Im),
    .io_in_22_Re(PermutationModuleStreamed_io_in_22_Re),
    .io_in_22_Im(PermutationModuleStreamed_io_in_22_Im),
    .io_in_23_Re(PermutationModuleStreamed_io_in_23_Re),
    .io_in_23_Im(PermutationModuleStreamed_io_in_23_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_in_config_7(PermutationModuleStreamed_io_in_config_7),
    .io_in_config_8(PermutationModuleStreamed_io_in_config_8),
    .io_in_config_9(PermutationModuleStreamed_io_in_config_9),
    .io_in_config_10(PermutationModuleStreamed_io_in_config_10),
    .io_in_config_11(PermutationModuleStreamed_io_in_config_11),
    .io_in_config_12(PermutationModuleStreamed_io_in_config_12),
    .io_in_config_13(PermutationModuleStreamed_io_in_config_13),
    .io_in_config_14(PermutationModuleStreamed_io_in_config_14),
    .io_in_config_15(PermutationModuleStreamed_io_in_config_15),
    .io_in_config_16(PermutationModuleStreamed_io_in_config_16),
    .io_in_config_17(PermutationModuleStreamed_io_in_config_17),
    .io_in_config_18(PermutationModuleStreamed_io_in_config_18),
    .io_in_config_19(PermutationModuleStreamed_io_in_config_19),
    .io_in_config_20(PermutationModuleStreamed_io_in_config_20),
    .io_in_config_21(PermutationModuleStreamed_io_in_config_21),
    .io_in_config_22(PermutationModuleStreamed_io_in_config_22),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im),
    .io_out_8_Re(PermutationModuleStreamed_io_out_8_Re),
    .io_out_8_Im(PermutationModuleStreamed_io_out_8_Im),
    .io_out_9_Re(PermutationModuleStreamed_io_out_9_Re),
    .io_out_9_Im(PermutationModuleStreamed_io_out_9_Im),
    .io_out_10_Re(PermutationModuleStreamed_io_out_10_Re),
    .io_out_10_Im(PermutationModuleStreamed_io_out_10_Im),
    .io_out_11_Re(PermutationModuleStreamed_io_out_11_Re),
    .io_out_11_Im(PermutationModuleStreamed_io_out_11_Im),
    .io_out_12_Re(PermutationModuleStreamed_io_out_12_Re),
    .io_out_12_Im(PermutationModuleStreamed_io_out_12_Im),
    .io_out_13_Re(PermutationModuleStreamed_io_out_13_Re),
    .io_out_13_Im(PermutationModuleStreamed_io_out_13_Im),
    .io_out_14_Re(PermutationModuleStreamed_io_out_14_Re),
    .io_out_14_Im(PermutationModuleStreamed_io_out_14_Im),
    .io_out_15_Re(PermutationModuleStreamed_io_out_15_Re),
    .io_out_15_Im(PermutationModuleStreamed_io_out_15_Im),
    .io_out_16_Re(PermutationModuleStreamed_io_out_16_Re),
    .io_out_16_Im(PermutationModuleStreamed_io_out_16_Im),
    .io_out_17_Re(PermutationModuleStreamed_io_out_17_Re),
    .io_out_17_Im(PermutationModuleStreamed_io_out_17_Im),
    .io_out_18_Re(PermutationModuleStreamed_io_out_18_Re),
    .io_out_18_Im(PermutationModuleStreamed_io_out_18_Im),
    .io_out_19_Re(PermutationModuleStreamed_io_out_19_Re),
    .io_out_19_Im(PermutationModuleStreamed_io_out_19_Im),
    .io_out_20_Re(PermutationModuleStreamed_io_out_20_Re),
    .io_out_20_Im(PermutationModuleStreamed_io_out_20_Im),
    .io_out_21_Re(PermutationModuleStreamed_io_out_21_Re),
    .io_out_21_Im(PermutationModuleStreamed_io_out_21_Im),
    .io_out_22_Re(PermutationModuleStreamed_io_out_22_Re),
    .io_out_22_Im(PermutationModuleStreamed_io_out_22_Im),
    .io_out_23_Re(PermutationModuleStreamed_io_out_23_Re),
    .io_out_23_Im(PermutationModuleStreamed_io_out_23_Im)
  );
  M0_Config_ROM_7 M0_Config_ROM ( // @[FFTDesigns.scala 2751:29]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7),
    .io_out_8(M0_Config_ROM_io_out_8),
    .io_out_9(M0_Config_ROM_io_out_9),
    .io_out_10(M0_Config_ROM_io_out_10),
    .io_out_11(M0_Config_ROM_io_out_11),
    .io_out_12(M0_Config_ROM_io_out_12),
    .io_out_13(M0_Config_ROM_io_out_13),
    .io_out_14(M0_Config_ROM_io_out_14),
    .io_out_15(M0_Config_ROM_io_out_15),
    .io_out_16(M0_Config_ROM_io_out_16),
    .io_out_17(M0_Config_ROM_io_out_17),
    .io_out_18(M0_Config_ROM_io_out_18),
    .io_out_19(M0_Config_ROM_io_out_19),
    .io_out_20(M0_Config_ROM_io_out_20),
    .io_out_21(M0_Config_ROM_io_out_21),
    .io_out_22(M0_Config_ROM_io_out_22),
    .io_out_23(M0_Config_ROM_io_out_23)
  );
  M1_Config_ROM_7 M1_Config_ROM ( // @[FFTDesigns.scala 2752:29]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7),
    .io_out_8(M1_Config_ROM_io_out_8),
    .io_out_9(M1_Config_ROM_io_out_9),
    .io_out_10(M1_Config_ROM_io_out_10),
    .io_out_11(M1_Config_ROM_io_out_11),
    .io_out_12(M1_Config_ROM_io_out_12),
    .io_out_13(M1_Config_ROM_io_out_13),
    .io_out_14(M1_Config_ROM_io_out_14),
    .io_out_15(M1_Config_ROM_io_out_15),
    .io_out_16(M1_Config_ROM_io_out_16),
    .io_out_17(M1_Config_ROM_io_out_17),
    .io_out_18(M1_Config_ROM_io_out_18),
    .io_out_19(M1_Config_ROM_io_out_19),
    .io_out_20(M1_Config_ROM_io_out_20),
    .io_out_21(M1_Config_ROM_io_out_21),
    .io_out_22(M1_Config_ROM_io_out_22),
    .io_out_23(M1_Config_ROM_io_out_23)
  );
  Streaming_Permute_Config_7 Streaming_Permute_Config ( // @[FFTDesigns.scala 2753:31]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6),
    .io_out_7(Streaming_Permute_Config_io_out_7),
    .io_out_8(Streaming_Permute_Config_io_out_8),
    .io_out_9(Streaming_Permute_Config_io_out_9),
    .io_out_10(Streaming_Permute_Config_io_out_10),
    .io_out_11(Streaming_Permute_Config_io_out_11),
    .io_out_12(Streaming_Permute_Config_io_out_12),
    .io_out_13(Streaming_Permute_Config_io_out_13),
    .io_out_14(Streaming_Permute_Config_io_out_14),
    .io_out_15(Streaming_Permute_Config_io_out_15),
    .io_out_16(Streaming_Permute_Config_io_out_16),
    .io_out_17(Streaming_Permute_Config_io_out_17),
    .io_out_18(Streaming_Permute_Config_io_out_18),
    .io_out_19(Streaming_Permute_Config_io_out_19),
    .io_out_20(Streaming_Permute_Config_io_out_20),
    .io_out_21(Streaming_Permute_Config_io_out_21),
    .io_out_22(Streaming_Permute_Config_io_out_22)
  );
  assign io_out_0_Re = RAM_Block_24_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_0_Im = RAM_Block_24_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_1_Re = RAM_Block_25_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_1_Im = RAM_Block_25_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_2_Re = RAM_Block_26_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_2_Im = RAM_Block_26_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_3_Re = RAM_Block_27_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_3_Im = RAM_Block_27_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_4_Re = RAM_Block_28_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_4_Im = RAM_Block_28_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_5_Re = RAM_Block_29_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_5_Im = RAM_Block_29_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_6_Re = RAM_Block_30_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_6_Im = RAM_Block_30_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_7_Re = RAM_Block_31_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_7_Im = RAM_Block_31_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_8_Re = RAM_Block_32_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_8_Im = RAM_Block_32_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_9_Re = RAM_Block_33_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_9_Im = RAM_Block_33_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_10_Re = RAM_Block_34_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_10_Im = RAM_Block_34_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_11_Re = RAM_Block_35_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_11_Im = RAM_Block_35_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_12_Re = RAM_Block_36_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_12_Im = RAM_Block_36_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_13_Re = RAM_Block_37_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_13_Im = RAM_Block_37_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_14_Re = RAM_Block_38_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_14_Im = RAM_Block_38_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_15_Re = RAM_Block_39_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_15_Im = RAM_Block_39_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_16_Re = RAM_Block_40_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_16_Im = RAM_Block_40_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_17_Re = RAM_Block_41_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_17_Im = RAM_Block_41_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_18_Re = RAM_Block_42_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_18_Im = RAM_Block_42_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_19_Re = RAM_Block_43_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_19_Im = RAM_Block_43_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_20_Re = RAM_Block_44_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_20_Im = RAM_Block_44_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_21_Re = RAM_Block_45_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_21_Im = RAM_Block_45_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_22_Re = RAM_Block_46_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_22_Im = RAM_Block_46_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_23_Re = RAM_Block_47_io_out_data_Re; // @[FFTDesigns.scala 2716:{23,23}]
  assign io_out_23_Im = RAM_Block_47_io_out_data_Im; // @[FFTDesigns.scala 2716:{23,23}]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = _GEN_2122[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_io_in_waddr = _GEN_2363[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_io_in_data_Re = M0_0_re ? _GEN_276 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_io_in_data_Im = M0_0_re ? _GEN_275 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_io_wr = M0_0_re & _GEN_273; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = _GEN_2132[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_1_io_in_waddr = _GEN_2368[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_1_io_in_data_Re = M0_0_re ? _GEN_356 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_1_io_in_data_Im = M0_0_re ? _GEN_355 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_1_io_wr = M0_0_re & _GEN_353; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = _GEN_2142[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_2_io_in_waddr = _GEN_2373[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_2_io_in_data_Re = M0_0_re ? _GEN_436 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_2_io_in_data_Im = M0_0_re ? _GEN_435 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_2_io_wr = M0_0_re & _GEN_433; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = _GEN_2152[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_3_io_in_waddr = _GEN_2378[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_3_io_in_data_Re = M0_0_re ? _GEN_516 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_3_io_in_data_Im = M0_0_re ? _GEN_515 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_3_io_wr = M0_0_re & _GEN_513; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = _GEN_2162[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_4_io_in_waddr = _GEN_2383[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_4_io_in_data_Re = M0_0_re ? _GEN_596 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_4_io_in_data_Im = M0_0_re ? _GEN_595 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_4_io_wr = M0_0_re & _GEN_593; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = _GEN_2172[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_5_io_in_waddr = _GEN_2388[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_5_io_in_data_Re = M0_0_re ? _GEN_676 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_5_io_in_data_Im = M0_0_re ? _GEN_675 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_5_io_wr = M0_0_re & _GEN_673; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = _GEN_2182[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_6_io_in_waddr = _GEN_2393[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_6_io_in_data_Re = M0_0_re ? _GEN_756 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_6_io_in_data_Im = M0_0_re ? _GEN_755 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_6_io_wr = M0_0_re & _GEN_753; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = _GEN_2192[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_7_io_in_waddr = _GEN_2398[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_7_io_in_data_Re = M0_0_re ? _GEN_836 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_7_io_in_data_Im = M0_0_re ? _GEN_835 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_7_io_wr = M0_0_re & _GEN_833; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = _GEN_2202[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_8_io_in_waddr = _GEN_2403[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_8_io_in_data_Re = M0_0_re ? _GEN_916 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_8_io_in_data_Im = M0_0_re ? _GEN_915 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_8_io_wr = M0_0_re & _GEN_913; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = _GEN_2212[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_9_io_in_waddr = _GEN_2408[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_9_io_in_data_Re = M0_0_re ? _GEN_996 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_9_io_in_data_Im = M0_0_re ? _GEN_995 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_9_io_wr = M0_0_re & _GEN_993; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = _GEN_2222[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_10_io_in_waddr = _GEN_2413[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_10_io_in_data_Re = M0_0_re ? _GEN_1076 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_10_io_in_data_Im = M0_0_re ? _GEN_1075 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_10_io_wr = M0_0_re & _GEN_1073; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = _GEN_2232[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_11_io_in_waddr = _GEN_2418[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_11_io_in_data_Re = M0_0_re ? _GEN_1156 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_11_io_in_data_Im = M0_0_re ? _GEN_1155 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_11_io_wr = M0_0_re & _GEN_1153; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = _GEN_2242[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_12_io_in_waddr = _GEN_2423[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_12_io_in_data_Re = M0_0_re ? _GEN_1236 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_12_io_in_data_Im = M0_0_re ? _GEN_1235 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_12_io_wr = M0_0_re & _GEN_1233; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = _GEN_2252[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_13_io_in_waddr = _GEN_2428[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_13_io_in_data_Re = M0_0_re ? _GEN_1316 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_13_io_in_data_Im = M0_0_re ? _GEN_1315 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_13_io_wr = M0_0_re & _GEN_1313; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = _GEN_2262[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_14_io_in_waddr = _GEN_2433[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_14_io_in_data_Re = M0_0_re ? _GEN_1396 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_14_io_in_data_Im = M0_0_re ? _GEN_1395 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_14_io_wr = M0_0_re & _GEN_1393; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = _GEN_2272[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_15_io_in_waddr = _GEN_2438[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_15_io_in_data_Re = M0_0_re ? _GEN_1476 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_15_io_in_data_Im = M0_0_re ? _GEN_1475 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_15_io_wr = M0_0_re & _GEN_1473; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_16_clock = clock;
  assign RAM_Block_16_io_in_raddr = _GEN_2282[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_16_io_in_waddr = _GEN_2443[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_16_io_in_data_Re = M0_0_re ? _GEN_1556 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_16_io_in_data_Im = M0_0_re ? _GEN_1555 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_16_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_16_io_wr = M0_0_re & _GEN_1553; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_16_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_17_clock = clock;
  assign RAM_Block_17_io_in_raddr = _GEN_2292[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_17_io_in_waddr = _GEN_2448[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_17_io_in_data_Re = M0_0_re ? _GEN_1636 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_17_io_in_data_Im = M0_0_re ? _GEN_1635 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_17_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_17_io_wr = M0_0_re & _GEN_1633; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_17_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_18_clock = clock;
  assign RAM_Block_18_io_in_raddr = _GEN_2302[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_18_io_in_waddr = _GEN_2453[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_18_io_in_data_Re = M0_0_re ? _GEN_1716 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_18_io_in_data_Im = M0_0_re ? _GEN_1715 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_18_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_18_io_wr = M0_0_re & _GEN_1713; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_18_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_19_clock = clock;
  assign RAM_Block_19_io_in_raddr = _GEN_2312[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_19_io_in_waddr = _GEN_2458[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_19_io_in_data_Re = M0_0_re ? _GEN_1796 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_19_io_in_data_Im = M0_0_re ? _GEN_1795 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_19_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_19_io_wr = M0_0_re & _GEN_1793; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_19_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_20_clock = clock;
  assign RAM_Block_20_io_in_raddr = _GEN_2322[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_20_io_in_waddr = _GEN_2463[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_20_io_in_data_Re = M0_0_re ? _GEN_1876 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_20_io_in_data_Im = M0_0_re ? _GEN_1875 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_20_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_20_io_wr = M0_0_re & _GEN_1873; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_20_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_21_clock = clock;
  assign RAM_Block_21_io_in_raddr = _GEN_2332[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_21_io_in_waddr = _GEN_2468[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_21_io_in_data_Re = M0_0_re ? _GEN_1956 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_21_io_in_data_Im = M0_0_re ? _GEN_1955 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_21_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_21_io_wr = M0_0_re & _GEN_1953; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_21_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_22_clock = clock;
  assign RAM_Block_22_io_in_raddr = _GEN_2342[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_22_io_in_waddr = _GEN_2473[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_22_io_in_data_Re = M0_0_re ? _GEN_2036 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_22_io_in_data_Im = M0_0_re ? _GEN_2035 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_22_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_22_io_wr = M0_0_re & _GEN_2033; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_22_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_23_clock = clock;
  assign RAM_Block_23_io_in_raddr = _GEN_2352[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_23_io_in_waddr = _GEN_2478[2:0]; // @[FFTDesigns.scala 2712:23]
  assign RAM_Block_23_io_in_data_Re = M0_0_re ? _GEN_2116 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_23_io_in_data_Im = M0_0_re ? _GEN_2115 : 32'h0; // @[FFTDesigns.scala 2757:33 2815:25]
  assign RAM_Block_23_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_23_io_wr = M0_0_re & _GEN_2113; // @[FFTDesigns.scala 2757:33 2809:20]
  assign RAM_Block_23_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_24_clock = clock;
  assign RAM_Block_24_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_24_io_in_waddr = _GEN_2124[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_24_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_24_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_24_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_24_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_24_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_25_clock = clock;
  assign RAM_Block_25_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_25_io_in_waddr = _GEN_2134[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_25_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_25_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_25_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_25_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_25_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_26_clock = clock;
  assign RAM_Block_26_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_26_io_in_waddr = _GEN_2144[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_26_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_26_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_26_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_26_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_26_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_27_clock = clock;
  assign RAM_Block_27_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_27_io_in_waddr = _GEN_2154[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_27_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_27_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_27_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_27_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_27_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_28_clock = clock;
  assign RAM_Block_28_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_28_io_in_waddr = _GEN_2164[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_28_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_28_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_28_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_28_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_28_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_29_clock = clock;
  assign RAM_Block_29_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_29_io_in_waddr = _GEN_2174[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_29_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_29_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_29_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_29_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_29_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_30_clock = clock;
  assign RAM_Block_30_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_30_io_in_waddr = _GEN_2184[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_30_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_30_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_30_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_30_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_30_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_31_clock = clock;
  assign RAM_Block_31_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_31_io_in_waddr = _GEN_2194[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_31_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_31_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_31_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_31_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_31_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_32_clock = clock;
  assign RAM_Block_32_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_32_io_in_waddr = _GEN_2204[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_32_io_in_data_Re = PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_32_io_in_data_Im = PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_32_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_32_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_32_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_33_clock = clock;
  assign RAM_Block_33_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_33_io_in_waddr = _GEN_2214[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_33_io_in_data_Re = PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_33_io_in_data_Im = PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_33_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_33_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_33_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_34_clock = clock;
  assign RAM_Block_34_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_34_io_in_waddr = _GEN_2224[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_34_io_in_data_Re = PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_34_io_in_data_Im = PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_34_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_34_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_34_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_35_clock = clock;
  assign RAM_Block_35_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_35_io_in_waddr = _GEN_2234[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_35_io_in_data_Re = PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_35_io_in_data_Im = PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_35_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_35_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_35_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_36_clock = clock;
  assign RAM_Block_36_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_36_io_in_waddr = _GEN_2244[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_36_io_in_data_Re = PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_36_io_in_data_Im = PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_36_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_36_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_36_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_37_clock = clock;
  assign RAM_Block_37_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_37_io_in_waddr = _GEN_2254[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_37_io_in_data_Re = PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_37_io_in_data_Im = PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_37_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_37_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_37_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_38_clock = clock;
  assign RAM_Block_38_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_38_io_in_waddr = _GEN_2264[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_38_io_in_data_Re = PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_38_io_in_data_Im = PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_38_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_38_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_38_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_39_clock = clock;
  assign RAM_Block_39_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_39_io_in_waddr = _GEN_2274[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_39_io_in_data_Re = PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_39_io_in_data_Im = PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_39_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_39_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_39_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_40_clock = clock;
  assign RAM_Block_40_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_40_io_in_waddr = _GEN_2284[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_40_io_in_data_Re = PermutationModuleStreamed_io_out_16_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_40_io_in_data_Im = PermutationModuleStreamed_io_out_16_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_40_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_40_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_40_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_41_clock = clock;
  assign RAM_Block_41_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_41_io_in_waddr = _GEN_2294[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_41_io_in_data_Re = PermutationModuleStreamed_io_out_17_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_41_io_in_data_Im = PermutationModuleStreamed_io_out_17_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_41_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_41_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_41_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_42_clock = clock;
  assign RAM_Block_42_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_42_io_in_waddr = _GEN_2304[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_42_io_in_data_Re = PermutationModuleStreamed_io_out_18_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_42_io_in_data_Im = PermutationModuleStreamed_io_out_18_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_42_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_42_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_42_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_43_clock = clock;
  assign RAM_Block_43_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_43_io_in_waddr = _GEN_2314[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_43_io_in_data_Re = PermutationModuleStreamed_io_out_19_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_43_io_in_data_Im = PermutationModuleStreamed_io_out_19_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_43_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_43_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_43_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_44_clock = clock;
  assign RAM_Block_44_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_44_io_in_waddr = _GEN_2324[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_44_io_in_data_Re = PermutationModuleStreamed_io_out_20_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_44_io_in_data_Im = PermutationModuleStreamed_io_out_20_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_44_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_44_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_44_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_45_clock = clock;
  assign RAM_Block_45_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_45_io_in_waddr = _GEN_2334[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_45_io_in_data_Re = PermutationModuleStreamed_io_out_21_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_45_io_in_data_Im = PermutationModuleStreamed_io_out_21_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_45_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_45_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_45_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_46_clock = clock;
  assign RAM_Block_46_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_46_io_in_waddr = _GEN_2344[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_46_io_in_data_Re = PermutationModuleStreamed_io_out_22_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_46_io_in_data_Im = PermutationModuleStreamed_io_out_22_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_46_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_46_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_46_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_47_clock = clock;
  assign RAM_Block_47_io_in_raddr = _GEN_2123[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_47_io_in_waddr = _GEN_2354[2:0]; // @[FFTDesigns.scala 2716:23]
  assign RAM_Block_47_io_in_data_Re = PermutationModuleStreamed_io_out_23_Re; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_47_io_in_data_Im = PermutationModuleStreamed_io_out_23_Im; // @[FFTDesigns.scala 2757:33 2783:25 2818:25]
  assign RAM_Block_47_io_re = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_47_io_wr = |_T; // @[FFTDesigns.scala 2757:28]
  assign RAM_Block_47_io_en = |_T; // @[FFTDesigns.scala 2757:28]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_8_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_8_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_9_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_9_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_10_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_10_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_11_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_11_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_12_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_12_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_13_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_13_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_14_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_14_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_15_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_15_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_16_Re = RAM_Block_16_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_16_Im = RAM_Block_16_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_17_Re = RAM_Block_17_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_17_Im = RAM_Block_17_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_18_Re = RAM_Block_18_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_18_Im = RAM_Block_18_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_19_Re = RAM_Block_19_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_19_Im = RAM_Block_19_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_20_Re = RAM_Block_20_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_20_Im = RAM_Block_20_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_21_Re = RAM_Block_21_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_21_Im = RAM_Block_21_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_22_Re = RAM_Block_22_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_22_Im = RAM_Block_22_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_23_Re = RAM_Block_23_io_out_data_Re; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_23_Im = RAM_Block_23_io_out_data_Im; // @[FFTDesigns.scala 2712:{23,23}]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_7 = Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_8 = Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_9 = Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_10 = Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_11 = Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_12 = Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_13 = Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_14 = Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_15 = Streaming_Permute_Config_io_out_15; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_16 = Streaming_Permute_Config_io_out_16; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_17 = Streaming_Permute_Config_io_out_17; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_18 = Streaming_Permute_Config_io_out_18; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_19 = Streaming_Permute_Config_io_out_19; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_20 = Streaming_Permute_Config_io_out_20; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_21 = Streaming_Permute_Config_io_out_21; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign PermutationModuleStreamed_io_in_config_22 = Streaming_Permute_Config_io_out_22; // @[FFTDesigns.scala 2757:33 2784:33 2819:33]
  assign M0_Config_ROM_io_in_cnt = cnt2; // @[FFTDesigns.scala 2829:24]
  assign M1_Config_ROM_io_in_cnt = cnt2; // @[FFTDesigns.scala 2830:24]
  assign Streaming_Permute_Config_io_in_cnt = cnt2; // @[FFTDesigns.scala 2831:26]
  always @(posedge clock) begin
    offset_switch <= M0_0_re & _GEN_5; // @[FFTDesigns.scala 2757:33 2825:23]
    if (reset) begin // @[FFTDesigns.scala 2755:25]
      cnt2 <= 2'h0; // @[FFTDesigns.scala 2755:25]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2757:33]
      if (cnt2 == 2'h3 & cnt == 3'h5) begin // @[FFTDesigns.scala 2758:69]
        cnt2 <= 2'h0; // @[FFTDesigns.scala 2759:16]
      end else if (!(_T_2)) begin // @[FFTDesigns.scala 2762:46]
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2767:16]
      end
    end
    if (reset) begin // @[FFTDesigns.scala 2756:24]
      cnt <= 3'h0; // @[FFTDesigns.scala 2756:24]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2757:33]
      if (cnt2 == 2'h3 & cnt == 3'h5) begin // @[FFTDesigns.scala 2758:69]
        cnt <= 3'h0; // @[FFTDesigns.scala 2760:15]
      end else if (_T_2) begin // @[FFTDesigns.scala 2762:46]
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2764:15]
      end else begin
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2768:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt2 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  cnt = _RAND_2[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAM_Block_mw(
  input         clock,
  input  [3:0]  io_in_raddr,
  input  [3:0]  io_in_waddr_0,
  input  [3:0]  io_in_waddr_1,
  input  [31:0] io_in_data_0_Re,
  input  [31:0] io_in_data_0_Im,
  input  [31:0] io_in_data_1_Re,
  input  [31:0] io_in_data_1_Im,
  input         io_re,
  input         io_wr_0,
  input         io_wr_1,
  input         io_en,
  output [31:0] io_out_data_Re,
  output [31:0] io_out_data_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_0_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_0_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_1_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_1_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_2_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_2_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_3_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_3_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_4_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_4_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_5_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_5_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_6_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_6_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_7_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_7_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_8_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_8_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_9_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_9_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_10_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_10_Im; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_11_Re; // @[FFTDesigns.scala 3313:18]
  reg [31:0] mem_11_Im; // @[FFTDesigns.scala 3313:18]
  wire [31:0] _GEN_0 = 4'h0 == io_in_waddr_0 ? io_in_data_0_Im : mem_0_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_1 = 4'h1 == io_in_waddr_0 ? io_in_data_0_Im : mem_1_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_2 = 4'h2 == io_in_waddr_0 ? io_in_data_0_Im : mem_2_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_3 = 4'h3 == io_in_waddr_0 ? io_in_data_0_Im : mem_3_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_4 = 4'h4 == io_in_waddr_0 ? io_in_data_0_Im : mem_4_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_5 = 4'h5 == io_in_waddr_0 ? io_in_data_0_Im : mem_5_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_6 = 4'h6 == io_in_waddr_0 ? io_in_data_0_Im : mem_6_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_7 = 4'h7 == io_in_waddr_0 ? io_in_data_0_Im : mem_7_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_8 = 4'h8 == io_in_waddr_0 ? io_in_data_0_Im : mem_8_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_9 = 4'h9 == io_in_waddr_0 ? io_in_data_0_Im : mem_9_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_10 = 4'ha == io_in_waddr_0 ? io_in_data_0_Im : mem_10_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_11 = 4'hb == io_in_waddr_0 ? io_in_data_0_Im : mem_11_Im; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_12 = 4'h0 == io_in_waddr_0 ? io_in_data_0_Re : mem_0_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_13 = 4'h1 == io_in_waddr_0 ? io_in_data_0_Re : mem_1_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_14 = 4'h2 == io_in_waddr_0 ? io_in_data_0_Re : mem_2_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_15 = 4'h3 == io_in_waddr_0 ? io_in_data_0_Re : mem_3_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_16 = 4'h4 == io_in_waddr_0 ? io_in_data_0_Re : mem_4_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_17 = 4'h5 == io_in_waddr_0 ? io_in_data_0_Re : mem_5_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_18 = 4'h6 == io_in_waddr_0 ? io_in_data_0_Re : mem_6_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_19 = 4'h7 == io_in_waddr_0 ? io_in_data_0_Re : mem_7_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_20 = 4'h8 == io_in_waddr_0 ? io_in_data_0_Re : mem_8_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_21 = 4'h9 == io_in_waddr_0 ? io_in_data_0_Re : mem_9_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_22 = 4'ha == io_in_waddr_0 ? io_in_data_0_Re : mem_10_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_23 = 4'hb == io_in_waddr_0 ? io_in_data_0_Re : mem_11_Re; // @[FFTDesigns.scala 3313:18 3317:{31,31}]
  wire [31:0] _GEN_24 = io_wr_0 ? _GEN_0 : mem_0_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_25 = io_wr_0 ? _GEN_1 : mem_1_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_26 = io_wr_0 ? _GEN_2 : mem_2_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_27 = io_wr_0 ? _GEN_3 : mem_3_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_28 = io_wr_0 ? _GEN_4 : mem_4_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_29 = io_wr_0 ? _GEN_5 : mem_5_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_30 = io_wr_0 ? _GEN_6 : mem_6_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_31 = io_wr_0 ? _GEN_7 : mem_7_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_32 = io_wr_0 ? _GEN_8 : mem_8_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_33 = io_wr_0 ? _GEN_9 : mem_9_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_34 = io_wr_0 ? _GEN_10 : mem_10_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_35 = io_wr_0 ? _GEN_11 : mem_11_Im; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_36 = io_wr_0 ? _GEN_12 : mem_0_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_37 = io_wr_0 ? _GEN_13 : mem_1_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_38 = io_wr_0 ? _GEN_14 : mem_2_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_39 = io_wr_0 ? _GEN_15 : mem_3_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_40 = io_wr_0 ? _GEN_16 : mem_4_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_41 = io_wr_0 ? _GEN_17 : mem_5_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_42 = io_wr_0 ? _GEN_18 : mem_6_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_43 = io_wr_0 ? _GEN_19 : mem_7_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_44 = io_wr_0 ? _GEN_20 : mem_8_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_45 = io_wr_0 ? _GEN_21 : mem_9_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_46 = io_wr_0 ? _GEN_22 : mem_10_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_47 = io_wr_0 ? _GEN_23 : mem_11_Re; // @[FFTDesigns.scala 3313:18 3316:23]
  wire [31:0] _GEN_97 = 4'h1 == io_in_raddr ? mem_1_Im : mem_0_Im; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_98 = 4'h2 == io_in_raddr ? mem_2_Im : _GEN_97; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_99 = 4'h3 == io_in_raddr ? mem_3_Im : _GEN_98; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_100 = 4'h4 == io_in_raddr ? mem_4_Im : _GEN_99; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_101 = 4'h5 == io_in_raddr ? mem_5_Im : _GEN_100; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_102 = 4'h6 == io_in_raddr ? mem_6_Im : _GEN_101; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_103 = 4'h7 == io_in_raddr ? mem_7_Im : _GEN_102; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_104 = 4'h8 == io_in_raddr ? mem_8_Im : _GEN_103; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_105 = 4'h9 == io_in_raddr ? mem_9_Im : _GEN_104; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_106 = 4'ha == io_in_raddr ? mem_10_Im : _GEN_105; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_107 = 4'hb == io_in_raddr ? mem_11_Im : _GEN_106; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_109 = 4'h1 == io_in_raddr ? mem_1_Re : mem_0_Re; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_110 = 4'h2 == io_in_raddr ? mem_2_Re : _GEN_109; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_111 = 4'h3 == io_in_raddr ? mem_3_Re : _GEN_110; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_112 = 4'h4 == io_in_raddr ? mem_4_Re : _GEN_111; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_113 = 4'h5 == io_in_raddr ? mem_5_Re : _GEN_112; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_114 = 4'h6 == io_in_raddr ? mem_6_Re : _GEN_113; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_115 = 4'h7 == io_in_raddr ? mem_7_Re : _GEN_114; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_116 = 4'h8 == io_in_raddr ? mem_8_Re : _GEN_115; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_117 = 4'h9 == io_in_raddr ? mem_9_Re : _GEN_116; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_118 = 4'ha == io_in_raddr ? mem_10_Re : _GEN_117; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_119 = 4'hb == io_in_raddr ? mem_11_Re : _GEN_118; // @[FFTDesigns.scala 3321:{21,21}]
  wire [31:0] _GEN_120 = io_re ? _GEN_107 : 32'h0; // @[FFTDesigns.scala 3320:18 3321:21 3324:24]
  wire [31:0] _GEN_121 = io_re ? _GEN_119 : 32'h0; // @[FFTDesigns.scala 3320:18 3321:21 3323:24]
  assign io_out_data_Re = io_en ? _GEN_121 : 32'h0; // @[FFTDesigns.scala 3314:16 3327:22]
  assign io_out_data_Im = io_en ? _GEN_120 : 32'h0; // @[FFTDesigns.scala 3314:16 3328:22]
  always @(posedge clock) begin
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h0 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_0_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_0_Re <= _GEN_36;
        end
      end else begin
        mem_0_Re <= _GEN_36;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h0 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_0_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_0_Im <= _GEN_24;
        end
      end else begin
        mem_0_Im <= _GEN_24;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h1 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_1_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_1_Re <= _GEN_37;
        end
      end else begin
        mem_1_Re <= _GEN_37;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h1 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_1_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_1_Im <= _GEN_25;
        end
      end else begin
        mem_1_Im <= _GEN_25;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h2 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_2_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_2_Re <= _GEN_38;
        end
      end else begin
        mem_2_Re <= _GEN_38;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h2 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_2_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_2_Im <= _GEN_26;
        end
      end else begin
        mem_2_Im <= _GEN_26;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h3 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_3_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_3_Re <= _GEN_39;
        end
      end else begin
        mem_3_Re <= _GEN_39;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h3 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_3_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_3_Im <= _GEN_27;
        end
      end else begin
        mem_3_Im <= _GEN_27;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h4 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_4_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_4_Re <= _GEN_40;
        end
      end else begin
        mem_4_Re <= _GEN_40;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h4 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_4_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_4_Im <= _GEN_28;
        end
      end else begin
        mem_4_Im <= _GEN_28;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h5 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_5_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_5_Re <= _GEN_41;
        end
      end else begin
        mem_5_Re <= _GEN_41;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h5 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_5_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_5_Im <= _GEN_29;
        end
      end else begin
        mem_5_Im <= _GEN_29;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h6 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_6_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_6_Re <= _GEN_42;
        end
      end else begin
        mem_6_Re <= _GEN_42;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h6 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_6_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_6_Im <= _GEN_30;
        end
      end else begin
        mem_6_Im <= _GEN_30;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h7 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_7_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_7_Re <= _GEN_43;
        end
      end else begin
        mem_7_Re <= _GEN_43;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h7 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_7_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_7_Im <= _GEN_31;
        end
      end else begin
        mem_7_Im <= _GEN_31;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h8 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_8_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_8_Re <= _GEN_44;
        end
      end else begin
        mem_8_Re <= _GEN_44;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h8 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_8_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_8_Im <= _GEN_32;
        end
      end else begin
        mem_8_Im <= _GEN_32;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h9 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_9_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_9_Re <= _GEN_45;
        end
      end else begin
        mem_9_Re <= _GEN_45;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'h9 == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_9_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_9_Im <= _GEN_33;
        end
      end else begin
        mem_9_Im <= _GEN_33;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'ha == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_10_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_10_Re <= _GEN_46;
        end
      end else begin
        mem_10_Re <= _GEN_46;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'ha == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_10_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_10_Im <= _GEN_34;
        end
      end else begin
        mem_10_Im <= _GEN_34;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'hb == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_11_Re <= io_in_data_1_Re; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_11_Re <= _GEN_47;
        end
      end else begin
        mem_11_Re <= _GEN_47;
      end
    end
    if (io_en) begin // @[FFTDesigns.scala 3314:16]
      if (io_wr_1) begin // @[FFTDesigns.scala 3316:23]
        if (4'hb == io_in_waddr_1) begin // @[FFTDesigns.scala 3317:31]
          mem_11_Im <= io_in_data_1_Im; // @[FFTDesigns.scala 3317:31]
        end else begin
          mem_11_Im <= _GEN_35;
        end
      end else begin
        mem_11_Im <= _GEN_35;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_Re = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_Im = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_1_Re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mem_1_Im = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  mem_2_Re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mem_2_Im = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mem_3_Re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  mem_3_Im = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  mem_4_Re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  mem_4_Im = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  mem_5_Re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mem_5_Im = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mem_6_Re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  mem_6_Im = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  mem_7_Re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  mem_7_Im = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  mem_8_Re = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mem_8_Im = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mem_9_Re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mem_9_Im = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mem_10_Re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mem_10_Im = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_11_Re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mem_11_Im = _RAND_23[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PermutationsWithStreaming_mr_1(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  input         io_in_en_2,
  input         io_in_en_3,
  input         io_in_en_4,
  input         io_in_en_5,
  input         io_in_en_6,
  input         io_in_en_7,
  input         io_in_en_8,
  input         io_in_en_9,
  input         io_in_en_10,
  input         io_in_en_11,
  input         io_in_en_12,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  wire  RAM_Block_mw_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_1_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_1_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_1_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_1_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_1_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_2_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_2_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_2_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_2_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_2_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_3_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_3_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_3_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_3_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_3_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_4_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_4_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_4_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_4_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_4_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_5_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_5_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_5_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_5_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_5_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_6_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_6_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_6_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_6_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_6_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_7_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_7_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_7_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_7_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_7_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_8_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_8_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_8_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_8_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_8_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_8_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_8_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_8_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_8_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_8_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_8_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_8_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_8_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_8_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_9_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_9_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_9_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_9_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_9_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_9_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_9_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_9_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_9_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_9_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_9_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_9_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_9_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_9_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_10_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_10_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_10_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_10_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_10_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_10_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_10_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_10_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_10_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_10_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_10_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_10_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_10_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_10_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_11_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_11_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_11_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_11_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_11_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_11_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_11_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_11_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_11_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_11_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_11_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_11_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_11_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_11_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_12_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_12_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_12_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_12_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_12_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_12_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_12_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_12_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_12_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_12_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_12_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_12_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_12_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_12_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_13_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_13_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_13_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_13_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_13_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_13_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_13_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_13_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_13_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_13_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_13_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_13_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_13_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_13_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_14_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_14_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_14_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_14_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_14_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_14_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_14_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_14_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_14_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_14_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_14_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_14_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_14_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_14_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_15_clock; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_15_io_in_raddr; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_15_io_in_waddr_0; // @[FFTDesigns.scala 2837:26]
  wire [3:0] RAM_Block_mw_15_io_in_waddr_1; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_15_io_in_data_0_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_15_io_in_data_0_Im; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_15_io_in_data_1_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_15_io_in_data_1_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_15_io_re; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_15_io_wr_0; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_15_io_wr_1; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_mw_15_io_en; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_15_io_out_data_Re; // @[FFTDesigns.scala 2837:26]
  wire [31:0] RAM_Block_mw_15_io_out_data_Im; // @[FFTDesigns.scala 2837:26]
  wire  RAM_Block_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_1_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_1_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_1_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_1_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_1_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_1_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_1_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_1_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_2_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_2_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_2_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_2_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_2_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_2_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_2_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_2_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_3_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_3_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_3_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_3_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_3_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_3_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_3_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_3_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_4_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_4_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_4_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_4_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_4_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_4_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_4_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_4_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_5_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_5_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_5_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_5_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_5_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_5_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_5_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_5_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_6_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_6_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_6_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_6_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_6_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_6_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_6_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_6_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_7_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_7_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_7_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_7_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_7_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_7_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_7_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_7_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_8_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_8_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_8_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_8_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_8_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_8_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_8_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_8_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_9_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_9_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_9_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_9_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_9_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_9_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_9_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_9_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_10_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_10_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_10_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_10_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_10_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_10_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_10_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_10_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_11_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_11_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_11_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_11_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_11_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_11_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_11_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_11_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_12_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_12_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_12_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_12_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_12_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_12_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_12_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_12_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_13_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_13_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_13_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_13_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_13_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_13_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_13_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_13_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_14_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_14_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_14_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_14_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_14_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_14_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_14_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_14_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_15_clock; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_15_io_in_raddr; // @[FFTDesigns.scala 2841:26]
  wire [3:0] RAM_Block_15_io_in_waddr; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_15_io_in_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_15_io_in_data_Im; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_15_io_re; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_15_io_wr; // @[FFTDesigns.scala 2841:26]
  wire  RAM_Block_15_io_en; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2841:26]
  wire [31:0] RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2841:26]
  wire [31:0] PermutationModuleStreamed_io_in_0_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_0_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_1_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_1_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_2_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_2_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_3_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_3_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_4_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_4_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_5_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_5_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_6_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_6_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_7_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_7_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_8_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_8_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_9_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_9_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_10_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_10_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_11_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_11_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_12_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_12_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_13_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_13_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_14_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_14_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_15_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_in_15_Im; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_0; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_1; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_2; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_3; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_4; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_5; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_6; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_7; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_8; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_9; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_10; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_11; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_12; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_13; // @[FFTDesigns.scala 2907:28]
  wire [3:0] PermutationModuleStreamed_io_in_config_14; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2907:28]
  wire [31:0] PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2907:28]
  wire [2:0] M0_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_0; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_1; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_2; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_3; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_4; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_5; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_6; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_7; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_8; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_9; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_10; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_11; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_12; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_13; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_14; // @[FFTDesigns.scala 2908:29]
  wire [3:0] M0_Config_ROM_io_out_15; // @[FFTDesigns.scala 2908:29]
  wire [2:0] M1_Config_ROM_io_in_cnt; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_0; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_1; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_2; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_3; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_4; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_5; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_6; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_7; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_8; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_9; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_10; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_11; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_12; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_13; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_14; // @[FFTDesigns.scala 2909:29]
  wire [3:0] M1_Config_ROM_io_out_15; // @[FFTDesigns.scala 2909:29]
  wire [2:0] Streaming_Permute_Config_io_in_cnt; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2910:31]
  wire [3:0] Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2910:31]
  reg  offset_switch; // @[FFTDesigns.scala 2710:28]
  reg [31:0] input_delay_registers_0_0_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_0_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_1_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_1_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_2_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_2_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_3_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_3_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_4_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_4_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_5_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_5_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_6_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_6_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_7_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_7_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_8_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_8_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_9_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_9_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_10_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_10_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_11_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_11_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_12_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_12_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_13_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_13_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_14_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_14_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_15_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_15_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_16_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_16_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_17_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_17_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_18_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_18_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_19_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_19_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_20_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_20_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_21_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_21_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_22_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_22_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_23_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_0_23_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_1_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_1_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_2_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_2_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_3_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_3_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_4_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_4_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_5_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_5_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_6_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_6_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_7_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_7_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_8_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_8_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_9_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_9_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_10_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_10_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_11_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_11_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_12_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_12_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_13_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_13_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_14_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_14_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_15_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_15_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_16_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_16_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_17_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_17_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_18_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_18_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_19_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_19_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_20_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_20_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_21_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_21_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_22_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_22_Im; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_23_Re; // @[FFTDesigns.scala 2834:42]
  reg [31:0] input_delay_registers_1_23_Im; // @[FFTDesigns.scala 2834:42]
  reg [2:0] cnt2; // @[FFTDesigns.scala 2912:25]
  reg [1:0] cnt; // @[FFTDesigns.scala 2913:24]
  wire [5:0] lo = {io_in_en_5,io_in_en_4,io_in_en_3,io_in_en_2,io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2914:21]
  wire [12:0] _T = {io_in_en_12,io_in_en_11,io_in_en_10,io_in_en_9,io_in_en_8,io_in_en_7,io_in_en_6,lo}; // @[FFTDesigns.scala 2914:21]
  wire  M0_0_re = |_T; // @[FFTDesigns.scala 2914:28]
  wire  _T_3 = cnt == 2'h3; // @[FFTDesigns.scala 2922:46]
  wire  _offset_switch_T = ~offset_switch; // @[FFTDesigns.scala 2925:28]
  wire [2:0] _cnt2_T_1 = cnt2 + 3'h1; // @[FFTDesigns.scala 2928:24]
  wire [1:0] _cnt_T_1 = cnt + 2'h1; // @[FFTDesigns.scala 2933:24]
  wire [1:0] _GEN_0 = cnt2 >= 3'h2 ? _cnt_T_1 : 2'h0; // @[FFTDesigns.scala 2932:32 2933:17 2935:17]
  wire  _GEN_6 = cnt2 == 3'h5 & cnt == 2'h3 ? ~offset_switch : offset_switch; // @[FFTDesigns.scala 2922:69 2925:25]
  wire [3:0] _M0_0_in_raddr_T_1 = 3'h6 * _offset_switch_T; // @[FFTDesigns.scala 2950:56]
  wire [3:0] _M0_0_in_raddr_T_3 = M0_Config_ROM_io_out_0 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _GEN_2318 = {{1'd0}, cnt2}; // @[FFTDesigns.scala 2951:34]
  wire [3:0] _M1_0_in_raddr_T_3 = _GEN_2318 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2951:34]
  wire [3:0] _M1_0_in_waddr_T = 3'h6 * offset_switch; // @[FFTDesigns.scala 2952:56]
  wire [3:0] _M1_0_in_waddr_T_2 = M1_Config_ROM_io_out_0 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_1_in_raddr_T_3 = M0_Config_ROM_io_out_1 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_1_in_waddr_T_2 = M1_Config_ROM_io_out_1 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_2_in_raddr_T_3 = M0_Config_ROM_io_out_2 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_2_in_waddr_T_2 = M1_Config_ROM_io_out_2 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_3_in_raddr_T_3 = M0_Config_ROM_io_out_3 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_3_in_waddr_T_2 = M1_Config_ROM_io_out_3 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_4_in_raddr_T_3 = M0_Config_ROM_io_out_4 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_4_in_waddr_T_2 = M1_Config_ROM_io_out_4 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_5_in_raddr_T_3 = M0_Config_ROM_io_out_5 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_5_in_waddr_T_2 = M1_Config_ROM_io_out_5 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_6_in_raddr_T_3 = M0_Config_ROM_io_out_6 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_6_in_waddr_T_2 = M1_Config_ROM_io_out_6 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_7_in_raddr_T_3 = M0_Config_ROM_io_out_7 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_7_in_waddr_T_2 = M1_Config_ROM_io_out_7 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_8_in_raddr_T_3 = M0_Config_ROM_io_out_8 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_8_in_waddr_T_2 = M1_Config_ROM_io_out_8 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_9_in_raddr_T_3 = M0_Config_ROM_io_out_9 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_9_in_waddr_T_2 = M1_Config_ROM_io_out_9 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_10_in_raddr_T_3 = M0_Config_ROM_io_out_10 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_10_in_waddr_T_2 = M1_Config_ROM_io_out_10 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_11_in_raddr_T_3 = M0_Config_ROM_io_out_11 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_11_in_waddr_T_2 = M1_Config_ROM_io_out_11 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_12_in_raddr_T_3 = M0_Config_ROM_io_out_12 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_12_in_waddr_T_2 = M1_Config_ROM_io_out_12 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_13_in_raddr_T_3 = M0_Config_ROM_io_out_13 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_13_in_waddr_T_2 = M1_Config_ROM_io_out_13 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_14_in_raddr_T_3 = M0_Config_ROM_io_out_14 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_14_in_waddr_T_2 = M1_Config_ROM_io_out_14 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [3:0] _M0_15_in_raddr_T_3 = M0_Config_ROM_io_out_15 + _M0_0_in_raddr_T_1; // @[FFTDesigns.scala 2950:46]
  wire [3:0] _M1_15_in_waddr_T_2 = M1_Config_ROM_io_out_15 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2952:46]
  wire [2:0] _GEN_12 = 2'h1 == cnt ? 3'h2 : 3'h0; // @[FFTDesigns.scala 2978:{55,55}]
  wire [2:0] _GEN_13 = 2'h2 == cnt ? 3'h3 : _GEN_12; // @[FFTDesigns.scala 2978:{55,55}]
  wire [2:0] _GEN_14 = 2'h3 == cnt ? 3'h5 : _GEN_13; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_2334 = {{1'd0}, _GEN_14}; // @[FFTDesigns.scala 2978:55]
  wire [3:0] _M0_0_in_waddr_0_T_2 = _GEN_2334 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2978:55]
  wire [4:0] _GEN_16 = 2'h1 == cnt ? 5'h8 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_17 = 2'h2 == cnt ? 5'h0 : _GEN_16; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_18 = 2'h3 == cnt ? 5'h8 : _GEN_17; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_20 = 5'h1 == _GEN_18 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_21 = 5'h2 == _GEN_18 ? input_delay_registers_1_2_Im : _GEN_20; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_22 = 5'h3 == _GEN_18 ? input_delay_registers_1_3_Im : _GEN_21; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_23 = 5'h4 == _GEN_18 ? input_delay_registers_1_4_Im : _GEN_22; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_24 = 5'h5 == _GEN_18 ? input_delay_registers_1_5_Im : _GEN_23; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_25 = 5'h6 == _GEN_18 ? input_delay_registers_1_6_Im : _GEN_24; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_26 = 5'h7 == _GEN_18 ? input_delay_registers_1_7_Im : _GEN_25; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_27 = 5'h8 == _GEN_18 ? input_delay_registers_1_8_Im : _GEN_26; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_28 = 5'h9 == _GEN_18 ? input_delay_registers_1_9_Im : _GEN_27; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_29 = 5'ha == _GEN_18 ? input_delay_registers_1_10_Im : _GEN_28; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_30 = 5'hb == _GEN_18 ? input_delay_registers_1_11_Im : _GEN_29; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_31 = 5'hc == _GEN_18 ? input_delay_registers_1_12_Im : _GEN_30; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_32 = 5'hd == _GEN_18 ? input_delay_registers_1_13_Im : _GEN_31; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_33 = 5'he == _GEN_18 ? input_delay_registers_1_14_Im : _GEN_32; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_34 = 5'hf == _GEN_18 ? input_delay_registers_1_15_Im : _GEN_33; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_35 = 5'h10 == _GEN_18 ? input_delay_registers_1_16_Im : _GEN_34; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_36 = 5'h11 == _GEN_18 ? input_delay_registers_1_17_Im : _GEN_35; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_37 = 5'h12 == _GEN_18 ? input_delay_registers_1_18_Im : _GEN_36; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_38 = 5'h13 == _GEN_18 ? input_delay_registers_1_19_Im : _GEN_37; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_39 = 5'h14 == _GEN_18 ? input_delay_registers_1_20_Im : _GEN_38; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_40 = 5'h15 == _GEN_18 ? input_delay_registers_1_21_Im : _GEN_39; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_41 = 5'h16 == _GEN_18 ? input_delay_registers_1_22_Im : _GEN_40; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_42 = 5'h17 == _GEN_18 ? input_delay_registers_1_23_Im : _GEN_41; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_44 = 5'h1 == _GEN_18 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_45 = 5'h2 == _GEN_18 ? input_delay_registers_1_2_Re : _GEN_44; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_46 = 5'h3 == _GEN_18 ? input_delay_registers_1_3_Re : _GEN_45; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_47 = 5'h4 == _GEN_18 ? input_delay_registers_1_4_Re : _GEN_46; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_48 = 5'h5 == _GEN_18 ? input_delay_registers_1_5_Re : _GEN_47; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_49 = 5'h6 == _GEN_18 ? input_delay_registers_1_6_Re : _GEN_48; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_50 = 5'h7 == _GEN_18 ? input_delay_registers_1_7_Re : _GEN_49; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_51 = 5'h8 == _GEN_18 ? input_delay_registers_1_8_Re : _GEN_50; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_52 = 5'h9 == _GEN_18 ? input_delay_registers_1_9_Re : _GEN_51; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_53 = 5'ha == _GEN_18 ? input_delay_registers_1_10_Re : _GEN_52; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_54 = 5'hb == _GEN_18 ? input_delay_registers_1_11_Re : _GEN_53; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_55 = 5'hc == _GEN_18 ? input_delay_registers_1_12_Re : _GEN_54; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_56 = 5'hd == _GEN_18 ? input_delay_registers_1_13_Re : _GEN_55; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_57 = 5'he == _GEN_18 ? input_delay_registers_1_14_Re : _GEN_56; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_58 = 5'hf == _GEN_18 ? input_delay_registers_1_15_Re : _GEN_57; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_59 = 5'h10 == _GEN_18 ? input_delay_registers_1_16_Re : _GEN_58; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_60 = 5'h11 == _GEN_18 ? input_delay_registers_1_17_Re : _GEN_59; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_61 = 5'h12 == _GEN_18 ? input_delay_registers_1_18_Re : _GEN_60; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_62 = 5'h13 == _GEN_18 ? input_delay_registers_1_19_Re : _GEN_61; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_63 = 5'h14 == _GEN_18 ? input_delay_registers_1_20_Re : _GEN_62; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_64 = 5'h15 == _GEN_18 ? input_delay_registers_1_21_Re : _GEN_63; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_65 = 5'h16 == _GEN_18 ? input_delay_registers_1_22_Re : _GEN_64; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_66 = 5'h17 == _GEN_18 ? input_delay_registers_1_23_Re : _GEN_65; // @[FFTDesigns.scala 2979:{32,32}]
  wire  _GEN_68 = 2'h1 == cnt ? 1'h0 : 1'h1; // @[FFTDesigns.scala 2977:{27,27}]
  wire  _GEN_70 = 2'h3 == cnt ? 1'h0 : 2'h2 == cnt | _GEN_68; // @[FFTDesigns.scala 2977:{27,27}]
  wire [2:0] _GEN_72 = 2'h1 == cnt ? 3'h0 : 3'h1; // @[FFTDesigns.scala 2978:{55,55}]
  wire [2:0] _GEN_73 = 2'h2 == cnt ? 3'h4 : _GEN_72; // @[FFTDesigns.scala 2978:{55,55}]
  wire [2:0] _GEN_74 = 2'h3 == cnt ? 3'h0 : _GEN_73; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_2336 = {{1'd0}, _GEN_74}; // @[FFTDesigns.scala 2978:55]
  wire [3:0] _M0_0_in_waddr_1_T_2 = _GEN_2336 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2978:55]
  wire [4:0] _GEN_76 = 2'h1 == cnt ? 5'h0 : 5'h10; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_77 = 2'h2 == cnt ? 5'h10 : _GEN_76; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_78 = 2'h3 == cnt ? 5'h0 : _GEN_77; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_80 = 5'h1 == _GEN_78 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_81 = 5'h2 == _GEN_78 ? input_delay_registers_1_2_Im : _GEN_80; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_82 = 5'h3 == _GEN_78 ? input_delay_registers_1_3_Im : _GEN_81; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_83 = 5'h4 == _GEN_78 ? input_delay_registers_1_4_Im : _GEN_82; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_84 = 5'h5 == _GEN_78 ? input_delay_registers_1_5_Im : _GEN_83; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_85 = 5'h6 == _GEN_78 ? input_delay_registers_1_6_Im : _GEN_84; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_86 = 5'h7 == _GEN_78 ? input_delay_registers_1_7_Im : _GEN_85; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_87 = 5'h8 == _GEN_78 ? input_delay_registers_1_8_Im : _GEN_86; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_88 = 5'h9 == _GEN_78 ? input_delay_registers_1_9_Im : _GEN_87; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_89 = 5'ha == _GEN_78 ? input_delay_registers_1_10_Im : _GEN_88; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_90 = 5'hb == _GEN_78 ? input_delay_registers_1_11_Im : _GEN_89; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_91 = 5'hc == _GEN_78 ? input_delay_registers_1_12_Im : _GEN_90; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_92 = 5'hd == _GEN_78 ? input_delay_registers_1_13_Im : _GEN_91; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_93 = 5'he == _GEN_78 ? input_delay_registers_1_14_Im : _GEN_92; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_94 = 5'hf == _GEN_78 ? input_delay_registers_1_15_Im : _GEN_93; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_95 = 5'h10 == _GEN_78 ? input_delay_registers_1_16_Im : _GEN_94; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_96 = 5'h11 == _GEN_78 ? input_delay_registers_1_17_Im : _GEN_95; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_97 = 5'h12 == _GEN_78 ? input_delay_registers_1_18_Im : _GEN_96; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_98 = 5'h13 == _GEN_78 ? input_delay_registers_1_19_Im : _GEN_97; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_99 = 5'h14 == _GEN_78 ? input_delay_registers_1_20_Im : _GEN_98; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_100 = 5'h15 == _GEN_78 ? input_delay_registers_1_21_Im : _GEN_99; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_101 = 5'h16 == _GEN_78 ? input_delay_registers_1_22_Im : _GEN_100; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_102 = 5'h17 == _GEN_78 ? input_delay_registers_1_23_Im : _GEN_101; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_104 = 5'h1 == _GEN_78 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_105 = 5'h2 == _GEN_78 ? input_delay_registers_1_2_Re : _GEN_104; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_106 = 5'h3 == _GEN_78 ? input_delay_registers_1_3_Re : _GEN_105; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_107 = 5'h4 == _GEN_78 ? input_delay_registers_1_4_Re : _GEN_106; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_108 = 5'h5 == _GEN_78 ? input_delay_registers_1_5_Re : _GEN_107; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_109 = 5'h6 == _GEN_78 ? input_delay_registers_1_6_Re : _GEN_108; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_110 = 5'h7 == _GEN_78 ? input_delay_registers_1_7_Re : _GEN_109; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_111 = 5'h8 == _GEN_78 ? input_delay_registers_1_8_Re : _GEN_110; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_112 = 5'h9 == _GEN_78 ? input_delay_registers_1_9_Re : _GEN_111; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_113 = 5'ha == _GEN_78 ? input_delay_registers_1_10_Re : _GEN_112; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_114 = 5'hb == _GEN_78 ? input_delay_registers_1_11_Re : _GEN_113; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_115 = 5'hc == _GEN_78 ? input_delay_registers_1_12_Re : _GEN_114; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_116 = 5'hd == _GEN_78 ? input_delay_registers_1_13_Re : _GEN_115; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_117 = 5'he == _GEN_78 ? input_delay_registers_1_14_Re : _GEN_116; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_118 = 5'hf == _GEN_78 ? input_delay_registers_1_15_Re : _GEN_117; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_119 = 5'h10 == _GEN_78 ? input_delay_registers_1_16_Re : _GEN_118; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_120 = 5'h11 == _GEN_78 ? input_delay_registers_1_17_Re : _GEN_119; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_121 = 5'h12 == _GEN_78 ? input_delay_registers_1_18_Re : _GEN_120; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_122 = 5'h13 == _GEN_78 ? input_delay_registers_1_19_Re : _GEN_121; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_123 = 5'h14 == _GEN_78 ? input_delay_registers_1_20_Re : _GEN_122; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_124 = 5'h15 == _GEN_78 ? input_delay_registers_1_21_Re : _GEN_123; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_125 = 5'h16 == _GEN_78 ? input_delay_registers_1_22_Re : _GEN_124; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_126 = 5'h17 == _GEN_78 ? input_delay_registers_1_23_Re : _GEN_125; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_136 = 2'h1 == cnt ? 5'h9 : 5'h1; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_137 = 2'h2 == cnt ? 5'h1 : _GEN_136; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_138 = 2'h3 == cnt ? 5'h9 : _GEN_137; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_140 = 5'h1 == _GEN_138 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_141 = 5'h2 == _GEN_138 ? input_delay_registers_1_2_Im : _GEN_140; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_142 = 5'h3 == _GEN_138 ? input_delay_registers_1_3_Im : _GEN_141; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_143 = 5'h4 == _GEN_138 ? input_delay_registers_1_4_Im : _GEN_142; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_144 = 5'h5 == _GEN_138 ? input_delay_registers_1_5_Im : _GEN_143; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_145 = 5'h6 == _GEN_138 ? input_delay_registers_1_6_Im : _GEN_144; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_146 = 5'h7 == _GEN_138 ? input_delay_registers_1_7_Im : _GEN_145; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_147 = 5'h8 == _GEN_138 ? input_delay_registers_1_8_Im : _GEN_146; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_148 = 5'h9 == _GEN_138 ? input_delay_registers_1_9_Im : _GEN_147; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_149 = 5'ha == _GEN_138 ? input_delay_registers_1_10_Im : _GEN_148; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_150 = 5'hb == _GEN_138 ? input_delay_registers_1_11_Im : _GEN_149; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_151 = 5'hc == _GEN_138 ? input_delay_registers_1_12_Im : _GEN_150; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_152 = 5'hd == _GEN_138 ? input_delay_registers_1_13_Im : _GEN_151; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_153 = 5'he == _GEN_138 ? input_delay_registers_1_14_Im : _GEN_152; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_154 = 5'hf == _GEN_138 ? input_delay_registers_1_15_Im : _GEN_153; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_155 = 5'h10 == _GEN_138 ? input_delay_registers_1_16_Im : _GEN_154; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_156 = 5'h11 == _GEN_138 ? input_delay_registers_1_17_Im : _GEN_155; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_157 = 5'h12 == _GEN_138 ? input_delay_registers_1_18_Im : _GEN_156; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_158 = 5'h13 == _GEN_138 ? input_delay_registers_1_19_Im : _GEN_157; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_159 = 5'h14 == _GEN_138 ? input_delay_registers_1_20_Im : _GEN_158; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_160 = 5'h15 == _GEN_138 ? input_delay_registers_1_21_Im : _GEN_159; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_161 = 5'h16 == _GEN_138 ? input_delay_registers_1_22_Im : _GEN_160; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_162 = 5'h17 == _GEN_138 ? input_delay_registers_1_23_Im : _GEN_161; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_164 = 5'h1 == _GEN_138 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_165 = 5'h2 == _GEN_138 ? input_delay_registers_1_2_Re : _GEN_164; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_166 = 5'h3 == _GEN_138 ? input_delay_registers_1_3_Re : _GEN_165; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_167 = 5'h4 == _GEN_138 ? input_delay_registers_1_4_Re : _GEN_166; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_168 = 5'h5 == _GEN_138 ? input_delay_registers_1_5_Re : _GEN_167; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_169 = 5'h6 == _GEN_138 ? input_delay_registers_1_6_Re : _GEN_168; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_170 = 5'h7 == _GEN_138 ? input_delay_registers_1_7_Re : _GEN_169; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_171 = 5'h8 == _GEN_138 ? input_delay_registers_1_8_Re : _GEN_170; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_172 = 5'h9 == _GEN_138 ? input_delay_registers_1_9_Re : _GEN_171; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_173 = 5'ha == _GEN_138 ? input_delay_registers_1_10_Re : _GEN_172; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_174 = 5'hb == _GEN_138 ? input_delay_registers_1_11_Re : _GEN_173; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_175 = 5'hc == _GEN_138 ? input_delay_registers_1_12_Re : _GEN_174; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_176 = 5'hd == _GEN_138 ? input_delay_registers_1_13_Re : _GEN_175; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_177 = 5'he == _GEN_138 ? input_delay_registers_1_14_Re : _GEN_176; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_178 = 5'hf == _GEN_138 ? input_delay_registers_1_15_Re : _GEN_177; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_179 = 5'h10 == _GEN_138 ? input_delay_registers_1_16_Re : _GEN_178; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_180 = 5'h11 == _GEN_138 ? input_delay_registers_1_17_Re : _GEN_179; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_181 = 5'h12 == _GEN_138 ? input_delay_registers_1_18_Re : _GEN_180; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_182 = 5'h13 == _GEN_138 ? input_delay_registers_1_19_Re : _GEN_181; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_183 = 5'h14 == _GEN_138 ? input_delay_registers_1_20_Re : _GEN_182; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_184 = 5'h15 == _GEN_138 ? input_delay_registers_1_21_Re : _GEN_183; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_185 = 5'h16 == _GEN_138 ? input_delay_registers_1_22_Re : _GEN_184; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_186 = 5'h17 == _GEN_138 ? input_delay_registers_1_23_Re : _GEN_185; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_196 = 2'h1 == cnt ? 5'h0 : 5'h11; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_197 = 2'h2 == cnt ? 5'h11 : _GEN_196; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_198 = 2'h3 == cnt ? 5'h0 : _GEN_197; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_200 = 5'h1 == _GEN_198 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_201 = 5'h2 == _GEN_198 ? input_delay_registers_1_2_Im : _GEN_200; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_202 = 5'h3 == _GEN_198 ? input_delay_registers_1_3_Im : _GEN_201; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_203 = 5'h4 == _GEN_198 ? input_delay_registers_1_4_Im : _GEN_202; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_204 = 5'h5 == _GEN_198 ? input_delay_registers_1_5_Im : _GEN_203; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_205 = 5'h6 == _GEN_198 ? input_delay_registers_1_6_Im : _GEN_204; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_206 = 5'h7 == _GEN_198 ? input_delay_registers_1_7_Im : _GEN_205; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_207 = 5'h8 == _GEN_198 ? input_delay_registers_1_8_Im : _GEN_206; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_208 = 5'h9 == _GEN_198 ? input_delay_registers_1_9_Im : _GEN_207; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_209 = 5'ha == _GEN_198 ? input_delay_registers_1_10_Im : _GEN_208; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_210 = 5'hb == _GEN_198 ? input_delay_registers_1_11_Im : _GEN_209; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_211 = 5'hc == _GEN_198 ? input_delay_registers_1_12_Im : _GEN_210; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_212 = 5'hd == _GEN_198 ? input_delay_registers_1_13_Im : _GEN_211; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_213 = 5'he == _GEN_198 ? input_delay_registers_1_14_Im : _GEN_212; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_214 = 5'hf == _GEN_198 ? input_delay_registers_1_15_Im : _GEN_213; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_215 = 5'h10 == _GEN_198 ? input_delay_registers_1_16_Im : _GEN_214; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_216 = 5'h11 == _GEN_198 ? input_delay_registers_1_17_Im : _GEN_215; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_217 = 5'h12 == _GEN_198 ? input_delay_registers_1_18_Im : _GEN_216; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_218 = 5'h13 == _GEN_198 ? input_delay_registers_1_19_Im : _GEN_217; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_219 = 5'h14 == _GEN_198 ? input_delay_registers_1_20_Im : _GEN_218; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_220 = 5'h15 == _GEN_198 ? input_delay_registers_1_21_Im : _GEN_219; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_221 = 5'h16 == _GEN_198 ? input_delay_registers_1_22_Im : _GEN_220; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_222 = 5'h17 == _GEN_198 ? input_delay_registers_1_23_Im : _GEN_221; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_224 = 5'h1 == _GEN_198 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_225 = 5'h2 == _GEN_198 ? input_delay_registers_1_2_Re : _GEN_224; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_226 = 5'h3 == _GEN_198 ? input_delay_registers_1_3_Re : _GEN_225; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_227 = 5'h4 == _GEN_198 ? input_delay_registers_1_4_Re : _GEN_226; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_228 = 5'h5 == _GEN_198 ? input_delay_registers_1_5_Re : _GEN_227; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_229 = 5'h6 == _GEN_198 ? input_delay_registers_1_6_Re : _GEN_228; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_230 = 5'h7 == _GEN_198 ? input_delay_registers_1_7_Re : _GEN_229; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_231 = 5'h8 == _GEN_198 ? input_delay_registers_1_8_Re : _GEN_230; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_232 = 5'h9 == _GEN_198 ? input_delay_registers_1_9_Re : _GEN_231; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_233 = 5'ha == _GEN_198 ? input_delay_registers_1_10_Re : _GEN_232; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_234 = 5'hb == _GEN_198 ? input_delay_registers_1_11_Re : _GEN_233; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_235 = 5'hc == _GEN_198 ? input_delay_registers_1_12_Re : _GEN_234; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_236 = 5'hd == _GEN_198 ? input_delay_registers_1_13_Re : _GEN_235; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_237 = 5'he == _GEN_198 ? input_delay_registers_1_14_Re : _GEN_236; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_238 = 5'hf == _GEN_198 ? input_delay_registers_1_15_Re : _GEN_237; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_239 = 5'h10 == _GEN_198 ? input_delay_registers_1_16_Re : _GEN_238; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_240 = 5'h11 == _GEN_198 ? input_delay_registers_1_17_Re : _GEN_239; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_241 = 5'h12 == _GEN_198 ? input_delay_registers_1_18_Re : _GEN_240; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_242 = 5'h13 == _GEN_198 ? input_delay_registers_1_19_Re : _GEN_241; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_243 = 5'h14 == _GEN_198 ? input_delay_registers_1_20_Re : _GEN_242; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_244 = 5'h15 == _GEN_198 ? input_delay_registers_1_21_Re : _GEN_243; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_245 = 5'h16 == _GEN_198 ? input_delay_registers_1_22_Re : _GEN_244; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_246 = 5'h17 == _GEN_198 ? input_delay_registers_1_23_Re : _GEN_245; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_256 = 2'h1 == cnt ? 5'ha : 5'h2; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_257 = 2'h2 == cnt ? 5'h2 : _GEN_256; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_258 = 2'h3 == cnt ? 5'ha : _GEN_257; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_260 = 5'h1 == _GEN_258 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_261 = 5'h2 == _GEN_258 ? input_delay_registers_1_2_Im : _GEN_260; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_262 = 5'h3 == _GEN_258 ? input_delay_registers_1_3_Im : _GEN_261; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_263 = 5'h4 == _GEN_258 ? input_delay_registers_1_4_Im : _GEN_262; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_264 = 5'h5 == _GEN_258 ? input_delay_registers_1_5_Im : _GEN_263; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_265 = 5'h6 == _GEN_258 ? input_delay_registers_1_6_Im : _GEN_264; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_266 = 5'h7 == _GEN_258 ? input_delay_registers_1_7_Im : _GEN_265; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_267 = 5'h8 == _GEN_258 ? input_delay_registers_1_8_Im : _GEN_266; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_268 = 5'h9 == _GEN_258 ? input_delay_registers_1_9_Im : _GEN_267; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_269 = 5'ha == _GEN_258 ? input_delay_registers_1_10_Im : _GEN_268; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_270 = 5'hb == _GEN_258 ? input_delay_registers_1_11_Im : _GEN_269; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_271 = 5'hc == _GEN_258 ? input_delay_registers_1_12_Im : _GEN_270; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_272 = 5'hd == _GEN_258 ? input_delay_registers_1_13_Im : _GEN_271; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_273 = 5'he == _GEN_258 ? input_delay_registers_1_14_Im : _GEN_272; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_274 = 5'hf == _GEN_258 ? input_delay_registers_1_15_Im : _GEN_273; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_275 = 5'h10 == _GEN_258 ? input_delay_registers_1_16_Im : _GEN_274; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_276 = 5'h11 == _GEN_258 ? input_delay_registers_1_17_Im : _GEN_275; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_277 = 5'h12 == _GEN_258 ? input_delay_registers_1_18_Im : _GEN_276; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_278 = 5'h13 == _GEN_258 ? input_delay_registers_1_19_Im : _GEN_277; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_279 = 5'h14 == _GEN_258 ? input_delay_registers_1_20_Im : _GEN_278; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_280 = 5'h15 == _GEN_258 ? input_delay_registers_1_21_Im : _GEN_279; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_281 = 5'h16 == _GEN_258 ? input_delay_registers_1_22_Im : _GEN_280; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_282 = 5'h17 == _GEN_258 ? input_delay_registers_1_23_Im : _GEN_281; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_284 = 5'h1 == _GEN_258 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_285 = 5'h2 == _GEN_258 ? input_delay_registers_1_2_Re : _GEN_284; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_286 = 5'h3 == _GEN_258 ? input_delay_registers_1_3_Re : _GEN_285; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_287 = 5'h4 == _GEN_258 ? input_delay_registers_1_4_Re : _GEN_286; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_288 = 5'h5 == _GEN_258 ? input_delay_registers_1_5_Re : _GEN_287; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_289 = 5'h6 == _GEN_258 ? input_delay_registers_1_6_Re : _GEN_288; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_290 = 5'h7 == _GEN_258 ? input_delay_registers_1_7_Re : _GEN_289; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_291 = 5'h8 == _GEN_258 ? input_delay_registers_1_8_Re : _GEN_290; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_292 = 5'h9 == _GEN_258 ? input_delay_registers_1_9_Re : _GEN_291; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_293 = 5'ha == _GEN_258 ? input_delay_registers_1_10_Re : _GEN_292; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_294 = 5'hb == _GEN_258 ? input_delay_registers_1_11_Re : _GEN_293; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_295 = 5'hc == _GEN_258 ? input_delay_registers_1_12_Re : _GEN_294; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_296 = 5'hd == _GEN_258 ? input_delay_registers_1_13_Re : _GEN_295; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_297 = 5'he == _GEN_258 ? input_delay_registers_1_14_Re : _GEN_296; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_298 = 5'hf == _GEN_258 ? input_delay_registers_1_15_Re : _GEN_297; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_299 = 5'h10 == _GEN_258 ? input_delay_registers_1_16_Re : _GEN_298; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_300 = 5'h11 == _GEN_258 ? input_delay_registers_1_17_Re : _GEN_299; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_301 = 5'h12 == _GEN_258 ? input_delay_registers_1_18_Re : _GEN_300; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_302 = 5'h13 == _GEN_258 ? input_delay_registers_1_19_Re : _GEN_301; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_303 = 5'h14 == _GEN_258 ? input_delay_registers_1_20_Re : _GEN_302; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_304 = 5'h15 == _GEN_258 ? input_delay_registers_1_21_Re : _GEN_303; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_305 = 5'h16 == _GEN_258 ? input_delay_registers_1_22_Re : _GEN_304; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_306 = 5'h17 == _GEN_258 ? input_delay_registers_1_23_Re : _GEN_305; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_316 = 2'h1 == cnt ? 5'h0 : 5'h12; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_317 = 2'h2 == cnt ? 5'h12 : _GEN_316; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_318 = 2'h3 == cnt ? 5'h0 : _GEN_317; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_320 = 5'h1 == _GEN_318 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_321 = 5'h2 == _GEN_318 ? input_delay_registers_1_2_Im : _GEN_320; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_322 = 5'h3 == _GEN_318 ? input_delay_registers_1_3_Im : _GEN_321; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_323 = 5'h4 == _GEN_318 ? input_delay_registers_1_4_Im : _GEN_322; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_324 = 5'h5 == _GEN_318 ? input_delay_registers_1_5_Im : _GEN_323; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_325 = 5'h6 == _GEN_318 ? input_delay_registers_1_6_Im : _GEN_324; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_326 = 5'h7 == _GEN_318 ? input_delay_registers_1_7_Im : _GEN_325; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_327 = 5'h8 == _GEN_318 ? input_delay_registers_1_8_Im : _GEN_326; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_328 = 5'h9 == _GEN_318 ? input_delay_registers_1_9_Im : _GEN_327; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_329 = 5'ha == _GEN_318 ? input_delay_registers_1_10_Im : _GEN_328; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_330 = 5'hb == _GEN_318 ? input_delay_registers_1_11_Im : _GEN_329; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_331 = 5'hc == _GEN_318 ? input_delay_registers_1_12_Im : _GEN_330; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_332 = 5'hd == _GEN_318 ? input_delay_registers_1_13_Im : _GEN_331; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_333 = 5'he == _GEN_318 ? input_delay_registers_1_14_Im : _GEN_332; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_334 = 5'hf == _GEN_318 ? input_delay_registers_1_15_Im : _GEN_333; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_335 = 5'h10 == _GEN_318 ? input_delay_registers_1_16_Im : _GEN_334; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_336 = 5'h11 == _GEN_318 ? input_delay_registers_1_17_Im : _GEN_335; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_337 = 5'h12 == _GEN_318 ? input_delay_registers_1_18_Im : _GEN_336; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_338 = 5'h13 == _GEN_318 ? input_delay_registers_1_19_Im : _GEN_337; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_339 = 5'h14 == _GEN_318 ? input_delay_registers_1_20_Im : _GEN_338; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_340 = 5'h15 == _GEN_318 ? input_delay_registers_1_21_Im : _GEN_339; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_341 = 5'h16 == _GEN_318 ? input_delay_registers_1_22_Im : _GEN_340; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_342 = 5'h17 == _GEN_318 ? input_delay_registers_1_23_Im : _GEN_341; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_344 = 5'h1 == _GEN_318 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_345 = 5'h2 == _GEN_318 ? input_delay_registers_1_2_Re : _GEN_344; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_346 = 5'h3 == _GEN_318 ? input_delay_registers_1_3_Re : _GEN_345; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_347 = 5'h4 == _GEN_318 ? input_delay_registers_1_4_Re : _GEN_346; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_348 = 5'h5 == _GEN_318 ? input_delay_registers_1_5_Re : _GEN_347; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_349 = 5'h6 == _GEN_318 ? input_delay_registers_1_6_Re : _GEN_348; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_350 = 5'h7 == _GEN_318 ? input_delay_registers_1_7_Re : _GEN_349; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_351 = 5'h8 == _GEN_318 ? input_delay_registers_1_8_Re : _GEN_350; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_352 = 5'h9 == _GEN_318 ? input_delay_registers_1_9_Re : _GEN_351; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_353 = 5'ha == _GEN_318 ? input_delay_registers_1_10_Re : _GEN_352; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_354 = 5'hb == _GEN_318 ? input_delay_registers_1_11_Re : _GEN_353; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_355 = 5'hc == _GEN_318 ? input_delay_registers_1_12_Re : _GEN_354; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_356 = 5'hd == _GEN_318 ? input_delay_registers_1_13_Re : _GEN_355; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_357 = 5'he == _GEN_318 ? input_delay_registers_1_14_Re : _GEN_356; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_358 = 5'hf == _GEN_318 ? input_delay_registers_1_15_Re : _GEN_357; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_359 = 5'h10 == _GEN_318 ? input_delay_registers_1_16_Re : _GEN_358; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_360 = 5'h11 == _GEN_318 ? input_delay_registers_1_17_Re : _GEN_359; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_361 = 5'h12 == _GEN_318 ? input_delay_registers_1_18_Re : _GEN_360; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_362 = 5'h13 == _GEN_318 ? input_delay_registers_1_19_Re : _GEN_361; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_363 = 5'h14 == _GEN_318 ? input_delay_registers_1_20_Re : _GEN_362; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_364 = 5'h15 == _GEN_318 ? input_delay_registers_1_21_Re : _GEN_363; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_365 = 5'h16 == _GEN_318 ? input_delay_registers_1_22_Re : _GEN_364; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_366 = 5'h17 == _GEN_318 ? input_delay_registers_1_23_Re : _GEN_365; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_376 = 2'h1 == cnt ? 5'hb : 5'h3; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_377 = 2'h2 == cnt ? 5'h3 : _GEN_376; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_378 = 2'h3 == cnt ? 5'hb : _GEN_377; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_380 = 5'h1 == _GEN_378 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_381 = 5'h2 == _GEN_378 ? input_delay_registers_1_2_Im : _GEN_380; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_382 = 5'h3 == _GEN_378 ? input_delay_registers_1_3_Im : _GEN_381; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_383 = 5'h4 == _GEN_378 ? input_delay_registers_1_4_Im : _GEN_382; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_384 = 5'h5 == _GEN_378 ? input_delay_registers_1_5_Im : _GEN_383; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_385 = 5'h6 == _GEN_378 ? input_delay_registers_1_6_Im : _GEN_384; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_386 = 5'h7 == _GEN_378 ? input_delay_registers_1_7_Im : _GEN_385; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_387 = 5'h8 == _GEN_378 ? input_delay_registers_1_8_Im : _GEN_386; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_388 = 5'h9 == _GEN_378 ? input_delay_registers_1_9_Im : _GEN_387; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_389 = 5'ha == _GEN_378 ? input_delay_registers_1_10_Im : _GEN_388; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_390 = 5'hb == _GEN_378 ? input_delay_registers_1_11_Im : _GEN_389; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_391 = 5'hc == _GEN_378 ? input_delay_registers_1_12_Im : _GEN_390; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_392 = 5'hd == _GEN_378 ? input_delay_registers_1_13_Im : _GEN_391; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_393 = 5'he == _GEN_378 ? input_delay_registers_1_14_Im : _GEN_392; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_394 = 5'hf == _GEN_378 ? input_delay_registers_1_15_Im : _GEN_393; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_395 = 5'h10 == _GEN_378 ? input_delay_registers_1_16_Im : _GEN_394; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_396 = 5'h11 == _GEN_378 ? input_delay_registers_1_17_Im : _GEN_395; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_397 = 5'h12 == _GEN_378 ? input_delay_registers_1_18_Im : _GEN_396; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_398 = 5'h13 == _GEN_378 ? input_delay_registers_1_19_Im : _GEN_397; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_399 = 5'h14 == _GEN_378 ? input_delay_registers_1_20_Im : _GEN_398; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_400 = 5'h15 == _GEN_378 ? input_delay_registers_1_21_Im : _GEN_399; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_401 = 5'h16 == _GEN_378 ? input_delay_registers_1_22_Im : _GEN_400; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_402 = 5'h17 == _GEN_378 ? input_delay_registers_1_23_Im : _GEN_401; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_404 = 5'h1 == _GEN_378 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_405 = 5'h2 == _GEN_378 ? input_delay_registers_1_2_Re : _GEN_404; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_406 = 5'h3 == _GEN_378 ? input_delay_registers_1_3_Re : _GEN_405; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_407 = 5'h4 == _GEN_378 ? input_delay_registers_1_4_Re : _GEN_406; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_408 = 5'h5 == _GEN_378 ? input_delay_registers_1_5_Re : _GEN_407; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_409 = 5'h6 == _GEN_378 ? input_delay_registers_1_6_Re : _GEN_408; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_410 = 5'h7 == _GEN_378 ? input_delay_registers_1_7_Re : _GEN_409; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_411 = 5'h8 == _GEN_378 ? input_delay_registers_1_8_Re : _GEN_410; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_412 = 5'h9 == _GEN_378 ? input_delay_registers_1_9_Re : _GEN_411; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_413 = 5'ha == _GEN_378 ? input_delay_registers_1_10_Re : _GEN_412; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_414 = 5'hb == _GEN_378 ? input_delay_registers_1_11_Re : _GEN_413; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_415 = 5'hc == _GEN_378 ? input_delay_registers_1_12_Re : _GEN_414; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_416 = 5'hd == _GEN_378 ? input_delay_registers_1_13_Re : _GEN_415; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_417 = 5'he == _GEN_378 ? input_delay_registers_1_14_Re : _GEN_416; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_418 = 5'hf == _GEN_378 ? input_delay_registers_1_15_Re : _GEN_417; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_419 = 5'h10 == _GEN_378 ? input_delay_registers_1_16_Re : _GEN_418; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_420 = 5'h11 == _GEN_378 ? input_delay_registers_1_17_Re : _GEN_419; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_421 = 5'h12 == _GEN_378 ? input_delay_registers_1_18_Re : _GEN_420; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_422 = 5'h13 == _GEN_378 ? input_delay_registers_1_19_Re : _GEN_421; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_423 = 5'h14 == _GEN_378 ? input_delay_registers_1_20_Re : _GEN_422; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_424 = 5'h15 == _GEN_378 ? input_delay_registers_1_21_Re : _GEN_423; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_425 = 5'h16 == _GEN_378 ? input_delay_registers_1_22_Re : _GEN_424; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_426 = 5'h17 == _GEN_378 ? input_delay_registers_1_23_Re : _GEN_425; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_436 = 2'h1 == cnt ? 5'h0 : 5'h13; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_437 = 2'h2 == cnt ? 5'h13 : _GEN_436; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_438 = 2'h3 == cnt ? 5'h0 : _GEN_437; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_440 = 5'h1 == _GEN_438 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_441 = 5'h2 == _GEN_438 ? input_delay_registers_1_2_Im : _GEN_440; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_442 = 5'h3 == _GEN_438 ? input_delay_registers_1_3_Im : _GEN_441; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_443 = 5'h4 == _GEN_438 ? input_delay_registers_1_4_Im : _GEN_442; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_444 = 5'h5 == _GEN_438 ? input_delay_registers_1_5_Im : _GEN_443; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_445 = 5'h6 == _GEN_438 ? input_delay_registers_1_6_Im : _GEN_444; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_446 = 5'h7 == _GEN_438 ? input_delay_registers_1_7_Im : _GEN_445; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_447 = 5'h8 == _GEN_438 ? input_delay_registers_1_8_Im : _GEN_446; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_448 = 5'h9 == _GEN_438 ? input_delay_registers_1_9_Im : _GEN_447; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_449 = 5'ha == _GEN_438 ? input_delay_registers_1_10_Im : _GEN_448; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_450 = 5'hb == _GEN_438 ? input_delay_registers_1_11_Im : _GEN_449; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_451 = 5'hc == _GEN_438 ? input_delay_registers_1_12_Im : _GEN_450; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_452 = 5'hd == _GEN_438 ? input_delay_registers_1_13_Im : _GEN_451; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_453 = 5'he == _GEN_438 ? input_delay_registers_1_14_Im : _GEN_452; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_454 = 5'hf == _GEN_438 ? input_delay_registers_1_15_Im : _GEN_453; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_455 = 5'h10 == _GEN_438 ? input_delay_registers_1_16_Im : _GEN_454; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_456 = 5'h11 == _GEN_438 ? input_delay_registers_1_17_Im : _GEN_455; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_457 = 5'h12 == _GEN_438 ? input_delay_registers_1_18_Im : _GEN_456; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_458 = 5'h13 == _GEN_438 ? input_delay_registers_1_19_Im : _GEN_457; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_459 = 5'h14 == _GEN_438 ? input_delay_registers_1_20_Im : _GEN_458; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_460 = 5'h15 == _GEN_438 ? input_delay_registers_1_21_Im : _GEN_459; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_461 = 5'h16 == _GEN_438 ? input_delay_registers_1_22_Im : _GEN_460; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_462 = 5'h17 == _GEN_438 ? input_delay_registers_1_23_Im : _GEN_461; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_464 = 5'h1 == _GEN_438 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_465 = 5'h2 == _GEN_438 ? input_delay_registers_1_2_Re : _GEN_464; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_466 = 5'h3 == _GEN_438 ? input_delay_registers_1_3_Re : _GEN_465; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_467 = 5'h4 == _GEN_438 ? input_delay_registers_1_4_Re : _GEN_466; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_468 = 5'h5 == _GEN_438 ? input_delay_registers_1_5_Re : _GEN_467; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_469 = 5'h6 == _GEN_438 ? input_delay_registers_1_6_Re : _GEN_468; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_470 = 5'h7 == _GEN_438 ? input_delay_registers_1_7_Re : _GEN_469; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_471 = 5'h8 == _GEN_438 ? input_delay_registers_1_8_Re : _GEN_470; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_472 = 5'h9 == _GEN_438 ? input_delay_registers_1_9_Re : _GEN_471; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_473 = 5'ha == _GEN_438 ? input_delay_registers_1_10_Re : _GEN_472; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_474 = 5'hb == _GEN_438 ? input_delay_registers_1_11_Re : _GEN_473; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_475 = 5'hc == _GEN_438 ? input_delay_registers_1_12_Re : _GEN_474; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_476 = 5'hd == _GEN_438 ? input_delay_registers_1_13_Re : _GEN_475; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_477 = 5'he == _GEN_438 ? input_delay_registers_1_14_Re : _GEN_476; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_478 = 5'hf == _GEN_438 ? input_delay_registers_1_15_Re : _GEN_477; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_479 = 5'h10 == _GEN_438 ? input_delay_registers_1_16_Re : _GEN_478; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_480 = 5'h11 == _GEN_438 ? input_delay_registers_1_17_Re : _GEN_479; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_481 = 5'h12 == _GEN_438 ? input_delay_registers_1_18_Re : _GEN_480; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_482 = 5'h13 == _GEN_438 ? input_delay_registers_1_19_Re : _GEN_481; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_483 = 5'h14 == _GEN_438 ? input_delay_registers_1_20_Re : _GEN_482; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_484 = 5'h15 == _GEN_438 ? input_delay_registers_1_21_Re : _GEN_483; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_485 = 5'h16 == _GEN_438 ? input_delay_registers_1_22_Re : _GEN_484; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_486 = 5'h17 == _GEN_438 ? input_delay_registers_1_23_Re : _GEN_485; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_496 = 2'h1 == cnt ? 5'hc : 5'h4; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_497 = 2'h2 == cnt ? 5'h4 : _GEN_496; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_498 = 2'h3 == cnt ? 5'hc : _GEN_497; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_500 = 5'h1 == _GEN_498 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_501 = 5'h2 == _GEN_498 ? input_delay_registers_1_2_Im : _GEN_500; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_502 = 5'h3 == _GEN_498 ? input_delay_registers_1_3_Im : _GEN_501; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_503 = 5'h4 == _GEN_498 ? input_delay_registers_1_4_Im : _GEN_502; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_504 = 5'h5 == _GEN_498 ? input_delay_registers_1_5_Im : _GEN_503; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_505 = 5'h6 == _GEN_498 ? input_delay_registers_1_6_Im : _GEN_504; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_506 = 5'h7 == _GEN_498 ? input_delay_registers_1_7_Im : _GEN_505; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_507 = 5'h8 == _GEN_498 ? input_delay_registers_1_8_Im : _GEN_506; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_508 = 5'h9 == _GEN_498 ? input_delay_registers_1_9_Im : _GEN_507; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_509 = 5'ha == _GEN_498 ? input_delay_registers_1_10_Im : _GEN_508; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_510 = 5'hb == _GEN_498 ? input_delay_registers_1_11_Im : _GEN_509; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_511 = 5'hc == _GEN_498 ? input_delay_registers_1_12_Im : _GEN_510; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_512 = 5'hd == _GEN_498 ? input_delay_registers_1_13_Im : _GEN_511; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_513 = 5'he == _GEN_498 ? input_delay_registers_1_14_Im : _GEN_512; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_514 = 5'hf == _GEN_498 ? input_delay_registers_1_15_Im : _GEN_513; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_515 = 5'h10 == _GEN_498 ? input_delay_registers_1_16_Im : _GEN_514; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_516 = 5'h11 == _GEN_498 ? input_delay_registers_1_17_Im : _GEN_515; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_517 = 5'h12 == _GEN_498 ? input_delay_registers_1_18_Im : _GEN_516; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_518 = 5'h13 == _GEN_498 ? input_delay_registers_1_19_Im : _GEN_517; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_519 = 5'h14 == _GEN_498 ? input_delay_registers_1_20_Im : _GEN_518; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_520 = 5'h15 == _GEN_498 ? input_delay_registers_1_21_Im : _GEN_519; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_521 = 5'h16 == _GEN_498 ? input_delay_registers_1_22_Im : _GEN_520; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_522 = 5'h17 == _GEN_498 ? input_delay_registers_1_23_Im : _GEN_521; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_524 = 5'h1 == _GEN_498 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_525 = 5'h2 == _GEN_498 ? input_delay_registers_1_2_Re : _GEN_524; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_526 = 5'h3 == _GEN_498 ? input_delay_registers_1_3_Re : _GEN_525; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_527 = 5'h4 == _GEN_498 ? input_delay_registers_1_4_Re : _GEN_526; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_528 = 5'h5 == _GEN_498 ? input_delay_registers_1_5_Re : _GEN_527; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_529 = 5'h6 == _GEN_498 ? input_delay_registers_1_6_Re : _GEN_528; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_530 = 5'h7 == _GEN_498 ? input_delay_registers_1_7_Re : _GEN_529; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_531 = 5'h8 == _GEN_498 ? input_delay_registers_1_8_Re : _GEN_530; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_532 = 5'h9 == _GEN_498 ? input_delay_registers_1_9_Re : _GEN_531; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_533 = 5'ha == _GEN_498 ? input_delay_registers_1_10_Re : _GEN_532; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_534 = 5'hb == _GEN_498 ? input_delay_registers_1_11_Re : _GEN_533; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_535 = 5'hc == _GEN_498 ? input_delay_registers_1_12_Re : _GEN_534; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_536 = 5'hd == _GEN_498 ? input_delay_registers_1_13_Re : _GEN_535; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_537 = 5'he == _GEN_498 ? input_delay_registers_1_14_Re : _GEN_536; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_538 = 5'hf == _GEN_498 ? input_delay_registers_1_15_Re : _GEN_537; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_539 = 5'h10 == _GEN_498 ? input_delay_registers_1_16_Re : _GEN_538; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_540 = 5'h11 == _GEN_498 ? input_delay_registers_1_17_Re : _GEN_539; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_541 = 5'h12 == _GEN_498 ? input_delay_registers_1_18_Re : _GEN_540; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_542 = 5'h13 == _GEN_498 ? input_delay_registers_1_19_Re : _GEN_541; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_543 = 5'h14 == _GEN_498 ? input_delay_registers_1_20_Re : _GEN_542; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_544 = 5'h15 == _GEN_498 ? input_delay_registers_1_21_Re : _GEN_543; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_545 = 5'h16 == _GEN_498 ? input_delay_registers_1_22_Re : _GEN_544; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_546 = 5'h17 == _GEN_498 ? input_delay_registers_1_23_Re : _GEN_545; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_556 = 2'h1 == cnt ? 5'h0 : 5'h14; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_557 = 2'h2 == cnt ? 5'h14 : _GEN_556; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_558 = 2'h3 == cnt ? 5'h0 : _GEN_557; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_560 = 5'h1 == _GEN_558 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_561 = 5'h2 == _GEN_558 ? input_delay_registers_1_2_Im : _GEN_560; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_562 = 5'h3 == _GEN_558 ? input_delay_registers_1_3_Im : _GEN_561; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_563 = 5'h4 == _GEN_558 ? input_delay_registers_1_4_Im : _GEN_562; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_564 = 5'h5 == _GEN_558 ? input_delay_registers_1_5_Im : _GEN_563; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_565 = 5'h6 == _GEN_558 ? input_delay_registers_1_6_Im : _GEN_564; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_566 = 5'h7 == _GEN_558 ? input_delay_registers_1_7_Im : _GEN_565; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_567 = 5'h8 == _GEN_558 ? input_delay_registers_1_8_Im : _GEN_566; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_568 = 5'h9 == _GEN_558 ? input_delay_registers_1_9_Im : _GEN_567; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_569 = 5'ha == _GEN_558 ? input_delay_registers_1_10_Im : _GEN_568; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_570 = 5'hb == _GEN_558 ? input_delay_registers_1_11_Im : _GEN_569; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_571 = 5'hc == _GEN_558 ? input_delay_registers_1_12_Im : _GEN_570; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_572 = 5'hd == _GEN_558 ? input_delay_registers_1_13_Im : _GEN_571; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_573 = 5'he == _GEN_558 ? input_delay_registers_1_14_Im : _GEN_572; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_574 = 5'hf == _GEN_558 ? input_delay_registers_1_15_Im : _GEN_573; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_575 = 5'h10 == _GEN_558 ? input_delay_registers_1_16_Im : _GEN_574; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_576 = 5'h11 == _GEN_558 ? input_delay_registers_1_17_Im : _GEN_575; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_577 = 5'h12 == _GEN_558 ? input_delay_registers_1_18_Im : _GEN_576; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_578 = 5'h13 == _GEN_558 ? input_delay_registers_1_19_Im : _GEN_577; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_579 = 5'h14 == _GEN_558 ? input_delay_registers_1_20_Im : _GEN_578; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_580 = 5'h15 == _GEN_558 ? input_delay_registers_1_21_Im : _GEN_579; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_581 = 5'h16 == _GEN_558 ? input_delay_registers_1_22_Im : _GEN_580; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_582 = 5'h17 == _GEN_558 ? input_delay_registers_1_23_Im : _GEN_581; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_584 = 5'h1 == _GEN_558 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_585 = 5'h2 == _GEN_558 ? input_delay_registers_1_2_Re : _GEN_584; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_586 = 5'h3 == _GEN_558 ? input_delay_registers_1_3_Re : _GEN_585; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_587 = 5'h4 == _GEN_558 ? input_delay_registers_1_4_Re : _GEN_586; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_588 = 5'h5 == _GEN_558 ? input_delay_registers_1_5_Re : _GEN_587; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_589 = 5'h6 == _GEN_558 ? input_delay_registers_1_6_Re : _GEN_588; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_590 = 5'h7 == _GEN_558 ? input_delay_registers_1_7_Re : _GEN_589; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_591 = 5'h8 == _GEN_558 ? input_delay_registers_1_8_Re : _GEN_590; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_592 = 5'h9 == _GEN_558 ? input_delay_registers_1_9_Re : _GEN_591; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_593 = 5'ha == _GEN_558 ? input_delay_registers_1_10_Re : _GEN_592; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_594 = 5'hb == _GEN_558 ? input_delay_registers_1_11_Re : _GEN_593; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_595 = 5'hc == _GEN_558 ? input_delay_registers_1_12_Re : _GEN_594; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_596 = 5'hd == _GEN_558 ? input_delay_registers_1_13_Re : _GEN_595; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_597 = 5'he == _GEN_558 ? input_delay_registers_1_14_Re : _GEN_596; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_598 = 5'hf == _GEN_558 ? input_delay_registers_1_15_Re : _GEN_597; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_599 = 5'h10 == _GEN_558 ? input_delay_registers_1_16_Re : _GEN_598; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_600 = 5'h11 == _GEN_558 ? input_delay_registers_1_17_Re : _GEN_599; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_601 = 5'h12 == _GEN_558 ? input_delay_registers_1_18_Re : _GEN_600; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_602 = 5'h13 == _GEN_558 ? input_delay_registers_1_19_Re : _GEN_601; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_603 = 5'h14 == _GEN_558 ? input_delay_registers_1_20_Re : _GEN_602; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_604 = 5'h15 == _GEN_558 ? input_delay_registers_1_21_Re : _GEN_603; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_605 = 5'h16 == _GEN_558 ? input_delay_registers_1_22_Re : _GEN_604; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_606 = 5'h17 == _GEN_558 ? input_delay_registers_1_23_Re : _GEN_605; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_616 = 2'h1 == cnt ? 5'hd : 5'h5; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_617 = 2'h2 == cnt ? 5'h5 : _GEN_616; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_618 = 2'h3 == cnt ? 5'hd : _GEN_617; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_620 = 5'h1 == _GEN_618 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_621 = 5'h2 == _GEN_618 ? input_delay_registers_1_2_Im : _GEN_620; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_622 = 5'h3 == _GEN_618 ? input_delay_registers_1_3_Im : _GEN_621; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_623 = 5'h4 == _GEN_618 ? input_delay_registers_1_4_Im : _GEN_622; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_624 = 5'h5 == _GEN_618 ? input_delay_registers_1_5_Im : _GEN_623; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_625 = 5'h6 == _GEN_618 ? input_delay_registers_1_6_Im : _GEN_624; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_626 = 5'h7 == _GEN_618 ? input_delay_registers_1_7_Im : _GEN_625; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_627 = 5'h8 == _GEN_618 ? input_delay_registers_1_8_Im : _GEN_626; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_628 = 5'h9 == _GEN_618 ? input_delay_registers_1_9_Im : _GEN_627; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_629 = 5'ha == _GEN_618 ? input_delay_registers_1_10_Im : _GEN_628; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_630 = 5'hb == _GEN_618 ? input_delay_registers_1_11_Im : _GEN_629; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_631 = 5'hc == _GEN_618 ? input_delay_registers_1_12_Im : _GEN_630; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_632 = 5'hd == _GEN_618 ? input_delay_registers_1_13_Im : _GEN_631; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_633 = 5'he == _GEN_618 ? input_delay_registers_1_14_Im : _GEN_632; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_634 = 5'hf == _GEN_618 ? input_delay_registers_1_15_Im : _GEN_633; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_635 = 5'h10 == _GEN_618 ? input_delay_registers_1_16_Im : _GEN_634; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_636 = 5'h11 == _GEN_618 ? input_delay_registers_1_17_Im : _GEN_635; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_637 = 5'h12 == _GEN_618 ? input_delay_registers_1_18_Im : _GEN_636; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_638 = 5'h13 == _GEN_618 ? input_delay_registers_1_19_Im : _GEN_637; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_639 = 5'h14 == _GEN_618 ? input_delay_registers_1_20_Im : _GEN_638; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_640 = 5'h15 == _GEN_618 ? input_delay_registers_1_21_Im : _GEN_639; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_641 = 5'h16 == _GEN_618 ? input_delay_registers_1_22_Im : _GEN_640; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_642 = 5'h17 == _GEN_618 ? input_delay_registers_1_23_Im : _GEN_641; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_644 = 5'h1 == _GEN_618 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_645 = 5'h2 == _GEN_618 ? input_delay_registers_1_2_Re : _GEN_644; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_646 = 5'h3 == _GEN_618 ? input_delay_registers_1_3_Re : _GEN_645; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_647 = 5'h4 == _GEN_618 ? input_delay_registers_1_4_Re : _GEN_646; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_648 = 5'h5 == _GEN_618 ? input_delay_registers_1_5_Re : _GEN_647; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_649 = 5'h6 == _GEN_618 ? input_delay_registers_1_6_Re : _GEN_648; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_650 = 5'h7 == _GEN_618 ? input_delay_registers_1_7_Re : _GEN_649; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_651 = 5'h8 == _GEN_618 ? input_delay_registers_1_8_Re : _GEN_650; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_652 = 5'h9 == _GEN_618 ? input_delay_registers_1_9_Re : _GEN_651; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_653 = 5'ha == _GEN_618 ? input_delay_registers_1_10_Re : _GEN_652; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_654 = 5'hb == _GEN_618 ? input_delay_registers_1_11_Re : _GEN_653; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_655 = 5'hc == _GEN_618 ? input_delay_registers_1_12_Re : _GEN_654; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_656 = 5'hd == _GEN_618 ? input_delay_registers_1_13_Re : _GEN_655; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_657 = 5'he == _GEN_618 ? input_delay_registers_1_14_Re : _GEN_656; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_658 = 5'hf == _GEN_618 ? input_delay_registers_1_15_Re : _GEN_657; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_659 = 5'h10 == _GEN_618 ? input_delay_registers_1_16_Re : _GEN_658; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_660 = 5'h11 == _GEN_618 ? input_delay_registers_1_17_Re : _GEN_659; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_661 = 5'h12 == _GEN_618 ? input_delay_registers_1_18_Re : _GEN_660; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_662 = 5'h13 == _GEN_618 ? input_delay_registers_1_19_Re : _GEN_661; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_663 = 5'h14 == _GEN_618 ? input_delay_registers_1_20_Re : _GEN_662; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_664 = 5'h15 == _GEN_618 ? input_delay_registers_1_21_Re : _GEN_663; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_665 = 5'h16 == _GEN_618 ? input_delay_registers_1_22_Re : _GEN_664; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_666 = 5'h17 == _GEN_618 ? input_delay_registers_1_23_Re : _GEN_665; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_676 = 2'h1 == cnt ? 5'h0 : 5'h15; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_677 = 2'h2 == cnt ? 5'h15 : _GEN_676; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_678 = 2'h3 == cnt ? 5'h0 : _GEN_677; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_680 = 5'h1 == _GEN_678 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_681 = 5'h2 == _GEN_678 ? input_delay_registers_1_2_Im : _GEN_680; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_682 = 5'h3 == _GEN_678 ? input_delay_registers_1_3_Im : _GEN_681; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_683 = 5'h4 == _GEN_678 ? input_delay_registers_1_4_Im : _GEN_682; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_684 = 5'h5 == _GEN_678 ? input_delay_registers_1_5_Im : _GEN_683; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_685 = 5'h6 == _GEN_678 ? input_delay_registers_1_6_Im : _GEN_684; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_686 = 5'h7 == _GEN_678 ? input_delay_registers_1_7_Im : _GEN_685; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_687 = 5'h8 == _GEN_678 ? input_delay_registers_1_8_Im : _GEN_686; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_688 = 5'h9 == _GEN_678 ? input_delay_registers_1_9_Im : _GEN_687; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_689 = 5'ha == _GEN_678 ? input_delay_registers_1_10_Im : _GEN_688; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_690 = 5'hb == _GEN_678 ? input_delay_registers_1_11_Im : _GEN_689; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_691 = 5'hc == _GEN_678 ? input_delay_registers_1_12_Im : _GEN_690; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_692 = 5'hd == _GEN_678 ? input_delay_registers_1_13_Im : _GEN_691; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_693 = 5'he == _GEN_678 ? input_delay_registers_1_14_Im : _GEN_692; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_694 = 5'hf == _GEN_678 ? input_delay_registers_1_15_Im : _GEN_693; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_695 = 5'h10 == _GEN_678 ? input_delay_registers_1_16_Im : _GEN_694; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_696 = 5'h11 == _GEN_678 ? input_delay_registers_1_17_Im : _GEN_695; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_697 = 5'h12 == _GEN_678 ? input_delay_registers_1_18_Im : _GEN_696; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_698 = 5'h13 == _GEN_678 ? input_delay_registers_1_19_Im : _GEN_697; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_699 = 5'h14 == _GEN_678 ? input_delay_registers_1_20_Im : _GEN_698; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_700 = 5'h15 == _GEN_678 ? input_delay_registers_1_21_Im : _GEN_699; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_701 = 5'h16 == _GEN_678 ? input_delay_registers_1_22_Im : _GEN_700; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_702 = 5'h17 == _GEN_678 ? input_delay_registers_1_23_Im : _GEN_701; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_704 = 5'h1 == _GEN_678 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_705 = 5'h2 == _GEN_678 ? input_delay_registers_1_2_Re : _GEN_704; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_706 = 5'h3 == _GEN_678 ? input_delay_registers_1_3_Re : _GEN_705; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_707 = 5'h4 == _GEN_678 ? input_delay_registers_1_4_Re : _GEN_706; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_708 = 5'h5 == _GEN_678 ? input_delay_registers_1_5_Re : _GEN_707; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_709 = 5'h6 == _GEN_678 ? input_delay_registers_1_6_Re : _GEN_708; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_710 = 5'h7 == _GEN_678 ? input_delay_registers_1_7_Re : _GEN_709; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_711 = 5'h8 == _GEN_678 ? input_delay_registers_1_8_Re : _GEN_710; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_712 = 5'h9 == _GEN_678 ? input_delay_registers_1_9_Re : _GEN_711; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_713 = 5'ha == _GEN_678 ? input_delay_registers_1_10_Re : _GEN_712; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_714 = 5'hb == _GEN_678 ? input_delay_registers_1_11_Re : _GEN_713; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_715 = 5'hc == _GEN_678 ? input_delay_registers_1_12_Re : _GEN_714; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_716 = 5'hd == _GEN_678 ? input_delay_registers_1_13_Re : _GEN_715; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_717 = 5'he == _GEN_678 ? input_delay_registers_1_14_Re : _GEN_716; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_718 = 5'hf == _GEN_678 ? input_delay_registers_1_15_Re : _GEN_717; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_719 = 5'h10 == _GEN_678 ? input_delay_registers_1_16_Re : _GEN_718; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_720 = 5'h11 == _GEN_678 ? input_delay_registers_1_17_Re : _GEN_719; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_721 = 5'h12 == _GEN_678 ? input_delay_registers_1_18_Re : _GEN_720; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_722 = 5'h13 == _GEN_678 ? input_delay_registers_1_19_Re : _GEN_721; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_723 = 5'h14 == _GEN_678 ? input_delay_registers_1_20_Re : _GEN_722; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_724 = 5'h15 == _GEN_678 ? input_delay_registers_1_21_Re : _GEN_723; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_725 = 5'h16 == _GEN_678 ? input_delay_registers_1_22_Re : _GEN_724; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_726 = 5'h17 == _GEN_678 ? input_delay_registers_1_23_Re : _GEN_725; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_736 = 2'h1 == cnt ? 5'he : 5'h6; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_737 = 2'h2 == cnt ? 5'h6 : _GEN_736; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_738 = 2'h3 == cnt ? 5'he : _GEN_737; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_740 = 5'h1 == _GEN_738 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_741 = 5'h2 == _GEN_738 ? input_delay_registers_1_2_Im : _GEN_740; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_742 = 5'h3 == _GEN_738 ? input_delay_registers_1_3_Im : _GEN_741; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_743 = 5'h4 == _GEN_738 ? input_delay_registers_1_4_Im : _GEN_742; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_744 = 5'h5 == _GEN_738 ? input_delay_registers_1_5_Im : _GEN_743; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_745 = 5'h6 == _GEN_738 ? input_delay_registers_1_6_Im : _GEN_744; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_746 = 5'h7 == _GEN_738 ? input_delay_registers_1_7_Im : _GEN_745; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_747 = 5'h8 == _GEN_738 ? input_delay_registers_1_8_Im : _GEN_746; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_748 = 5'h9 == _GEN_738 ? input_delay_registers_1_9_Im : _GEN_747; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_749 = 5'ha == _GEN_738 ? input_delay_registers_1_10_Im : _GEN_748; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_750 = 5'hb == _GEN_738 ? input_delay_registers_1_11_Im : _GEN_749; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_751 = 5'hc == _GEN_738 ? input_delay_registers_1_12_Im : _GEN_750; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_752 = 5'hd == _GEN_738 ? input_delay_registers_1_13_Im : _GEN_751; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_753 = 5'he == _GEN_738 ? input_delay_registers_1_14_Im : _GEN_752; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_754 = 5'hf == _GEN_738 ? input_delay_registers_1_15_Im : _GEN_753; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_755 = 5'h10 == _GEN_738 ? input_delay_registers_1_16_Im : _GEN_754; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_756 = 5'h11 == _GEN_738 ? input_delay_registers_1_17_Im : _GEN_755; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_757 = 5'h12 == _GEN_738 ? input_delay_registers_1_18_Im : _GEN_756; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_758 = 5'h13 == _GEN_738 ? input_delay_registers_1_19_Im : _GEN_757; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_759 = 5'h14 == _GEN_738 ? input_delay_registers_1_20_Im : _GEN_758; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_760 = 5'h15 == _GEN_738 ? input_delay_registers_1_21_Im : _GEN_759; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_761 = 5'h16 == _GEN_738 ? input_delay_registers_1_22_Im : _GEN_760; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_762 = 5'h17 == _GEN_738 ? input_delay_registers_1_23_Im : _GEN_761; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_764 = 5'h1 == _GEN_738 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_765 = 5'h2 == _GEN_738 ? input_delay_registers_1_2_Re : _GEN_764; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_766 = 5'h3 == _GEN_738 ? input_delay_registers_1_3_Re : _GEN_765; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_767 = 5'h4 == _GEN_738 ? input_delay_registers_1_4_Re : _GEN_766; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_768 = 5'h5 == _GEN_738 ? input_delay_registers_1_5_Re : _GEN_767; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_769 = 5'h6 == _GEN_738 ? input_delay_registers_1_6_Re : _GEN_768; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_770 = 5'h7 == _GEN_738 ? input_delay_registers_1_7_Re : _GEN_769; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_771 = 5'h8 == _GEN_738 ? input_delay_registers_1_8_Re : _GEN_770; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_772 = 5'h9 == _GEN_738 ? input_delay_registers_1_9_Re : _GEN_771; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_773 = 5'ha == _GEN_738 ? input_delay_registers_1_10_Re : _GEN_772; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_774 = 5'hb == _GEN_738 ? input_delay_registers_1_11_Re : _GEN_773; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_775 = 5'hc == _GEN_738 ? input_delay_registers_1_12_Re : _GEN_774; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_776 = 5'hd == _GEN_738 ? input_delay_registers_1_13_Re : _GEN_775; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_777 = 5'he == _GEN_738 ? input_delay_registers_1_14_Re : _GEN_776; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_778 = 5'hf == _GEN_738 ? input_delay_registers_1_15_Re : _GEN_777; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_779 = 5'h10 == _GEN_738 ? input_delay_registers_1_16_Re : _GEN_778; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_780 = 5'h11 == _GEN_738 ? input_delay_registers_1_17_Re : _GEN_779; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_781 = 5'h12 == _GEN_738 ? input_delay_registers_1_18_Re : _GEN_780; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_782 = 5'h13 == _GEN_738 ? input_delay_registers_1_19_Re : _GEN_781; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_783 = 5'h14 == _GEN_738 ? input_delay_registers_1_20_Re : _GEN_782; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_784 = 5'h15 == _GEN_738 ? input_delay_registers_1_21_Re : _GEN_783; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_785 = 5'h16 == _GEN_738 ? input_delay_registers_1_22_Re : _GEN_784; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_786 = 5'h17 == _GEN_738 ? input_delay_registers_1_23_Re : _GEN_785; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_796 = 2'h1 == cnt ? 5'h0 : 5'h16; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_797 = 2'h2 == cnt ? 5'h16 : _GEN_796; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_798 = 2'h3 == cnt ? 5'h0 : _GEN_797; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_800 = 5'h1 == _GEN_798 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_801 = 5'h2 == _GEN_798 ? input_delay_registers_1_2_Im : _GEN_800; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_802 = 5'h3 == _GEN_798 ? input_delay_registers_1_3_Im : _GEN_801; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_803 = 5'h4 == _GEN_798 ? input_delay_registers_1_4_Im : _GEN_802; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_804 = 5'h5 == _GEN_798 ? input_delay_registers_1_5_Im : _GEN_803; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_805 = 5'h6 == _GEN_798 ? input_delay_registers_1_6_Im : _GEN_804; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_806 = 5'h7 == _GEN_798 ? input_delay_registers_1_7_Im : _GEN_805; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_807 = 5'h8 == _GEN_798 ? input_delay_registers_1_8_Im : _GEN_806; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_808 = 5'h9 == _GEN_798 ? input_delay_registers_1_9_Im : _GEN_807; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_809 = 5'ha == _GEN_798 ? input_delay_registers_1_10_Im : _GEN_808; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_810 = 5'hb == _GEN_798 ? input_delay_registers_1_11_Im : _GEN_809; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_811 = 5'hc == _GEN_798 ? input_delay_registers_1_12_Im : _GEN_810; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_812 = 5'hd == _GEN_798 ? input_delay_registers_1_13_Im : _GEN_811; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_813 = 5'he == _GEN_798 ? input_delay_registers_1_14_Im : _GEN_812; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_814 = 5'hf == _GEN_798 ? input_delay_registers_1_15_Im : _GEN_813; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_815 = 5'h10 == _GEN_798 ? input_delay_registers_1_16_Im : _GEN_814; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_816 = 5'h11 == _GEN_798 ? input_delay_registers_1_17_Im : _GEN_815; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_817 = 5'h12 == _GEN_798 ? input_delay_registers_1_18_Im : _GEN_816; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_818 = 5'h13 == _GEN_798 ? input_delay_registers_1_19_Im : _GEN_817; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_819 = 5'h14 == _GEN_798 ? input_delay_registers_1_20_Im : _GEN_818; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_820 = 5'h15 == _GEN_798 ? input_delay_registers_1_21_Im : _GEN_819; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_821 = 5'h16 == _GEN_798 ? input_delay_registers_1_22_Im : _GEN_820; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_822 = 5'h17 == _GEN_798 ? input_delay_registers_1_23_Im : _GEN_821; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_824 = 5'h1 == _GEN_798 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_825 = 5'h2 == _GEN_798 ? input_delay_registers_1_2_Re : _GEN_824; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_826 = 5'h3 == _GEN_798 ? input_delay_registers_1_3_Re : _GEN_825; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_827 = 5'h4 == _GEN_798 ? input_delay_registers_1_4_Re : _GEN_826; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_828 = 5'h5 == _GEN_798 ? input_delay_registers_1_5_Re : _GEN_827; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_829 = 5'h6 == _GEN_798 ? input_delay_registers_1_6_Re : _GEN_828; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_830 = 5'h7 == _GEN_798 ? input_delay_registers_1_7_Re : _GEN_829; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_831 = 5'h8 == _GEN_798 ? input_delay_registers_1_8_Re : _GEN_830; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_832 = 5'h9 == _GEN_798 ? input_delay_registers_1_9_Re : _GEN_831; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_833 = 5'ha == _GEN_798 ? input_delay_registers_1_10_Re : _GEN_832; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_834 = 5'hb == _GEN_798 ? input_delay_registers_1_11_Re : _GEN_833; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_835 = 5'hc == _GEN_798 ? input_delay_registers_1_12_Re : _GEN_834; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_836 = 5'hd == _GEN_798 ? input_delay_registers_1_13_Re : _GEN_835; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_837 = 5'he == _GEN_798 ? input_delay_registers_1_14_Re : _GEN_836; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_838 = 5'hf == _GEN_798 ? input_delay_registers_1_15_Re : _GEN_837; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_839 = 5'h10 == _GEN_798 ? input_delay_registers_1_16_Re : _GEN_838; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_840 = 5'h11 == _GEN_798 ? input_delay_registers_1_17_Re : _GEN_839; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_841 = 5'h12 == _GEN_798 ? input_delay_registers_1_18_Re : _GEN_840; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_842 = 5'h13 == _GEN_798 ? input_delay_registers_1_19_Re : _GEN_841; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_843 = 5'h14 == _GEN_798 ? input_delay_registers_1_20_Re : _GEN_842; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_844 = 5'h15 == _GEN_798 ? input_delay_registers_1_21_Re : _GEN_843; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_845 = 5'h16 == _GEN_798 ? input_delay_registers_1_22_Re : _GEN_844; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_846 = 5'h17 == _GEN_798 ? input_delay_registers_1_23_Re : _GEN_845; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_856 = 2'h1 == cnt ? 5'hf : 5'h7; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_857 = 2'h2 == cnt ? 5'h7 : _GEN_856; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_858 = 2'h3 == cnt ? 5'hf : _GEN_857; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_860 = 5'h1 == _GEN_858 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_861 = 5'h2 == _GEN_858 ? input_delay_registers_1_2_Im : _GEN_860; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_862 = 5'h3 == _GEN_858 ? input_delay_registers_1_3_Im : _GEN_861; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_863 = 5'h4 == _GEN_858 ? input_delay_registers_1_4_Im : _GEN_862; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_864 = 5'h5 == _GEN_858 ? input_delay_registers_1_5_Im : _GEN_863; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_865 = 5'h6 == _GEN_858 ? input_delay_registers_1_6_Im : _GEN_864; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_866 = 5'h7 == _GEN_858 ? input_delay_registers_1_7_Im : _GEN_865; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_867 = 5'h8 == _GEN_858 ? input_delay_registers_1_8_Im : _GEN_866; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_868 = 5'h9 == _GEN_858 ? input_delay_registers_1_9_Im : _GEN_867; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_869 = 5'ha == _GEN_858 ? input_delay_registers_1_10_Im : _GEN_868; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_870 = 5'hb == _GEN_858 ? input_delay_registers_1_11_Im : _GEN_869; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_871 = 5'hc == _GEN_858 ? input_delay_registers_1_12_Im : _GEN_870; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_872 = 5'hd == _GEN_858 ? input_delay_registers_1_13_Im : _GEN_871; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_873 = 5'he == _GEN_858 ? input_delay_registers_1_14_Im : _GEN_872; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_874 = 5'hf == _GEN_858 ? input_delay_registers_1_15_Im : _GEN_873; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_875 = 5'h10 == _GEN_858 ? input_delay_registers_1_16_Im : _GEN_874; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_876 = 5'h11 == _GEN_858 ? input_delay_registers_1_17_Im : _GEN_875; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_877 = 5'h12 == _GEN_858 ? input_delay_registers_1_18_Im : _GEN_876; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_878 = 5'h13 == _GEN_858 ? input_delay_registers_1_19_Im : _GEN_877; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_879 = 5'h14 == _GEN_858 ? input_delay_registers_1_20_Im : _GEN_878; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_880 = 5'h15 == _GEN_858 ? input_delay_registers_1_21_Im : _GEN_879; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_881 = 5'h16 == _GEN_858 ? input_delay_registers_1_22_Im : _GEN_880; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_882 = 5'h17 == _GEN_858 ? input_delay_registers_1_23_Im : _GEN_881; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_884 = 5'h1 == _GEN_858 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_885 = 5'h2 == _GEN_858 ? input_delay_registers_1_2_Re : _GEN_884; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_886 = 5'h3 == _GEN_858 ? input_delay_registers_1_3_Re : _GEN_885; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_887 = 5'h4 == _GEN_858 ? input_delay_registers_1_4_Re : _GEN_886; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_888 = 5'h5 == _GEN_858 ? input_delay_registers_1_5_Re : _GEN_887; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_889 = 5'h6 == _GEN_858 ? input_delay_registers_1_6_Re : _GEN_888; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_890 = 5'h7 == _GEN_858 ? input_delay_registers_1_7_Re : _GEN_889; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_891 = 5'h8 == _GEN_858 ? input_delay_registers_1_8_Re : _GEN_890; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_892 = 5'h9 == _GEN_858 ? input_delay_registers_1_9_Re : _GEN_891; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_893 = 5'ha == _GEN_858 ? input_delay_registers_1_10_Re : _GEN_892; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_894 = 5'hb == _GEN_858 ? input_delay_registers_1_11_Re : _GEN_893; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_895 = 5'hc == _GEN_858 ? input_delay_registers_1_12_Re : _GEN_894; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_896 = 5'hd == _GEN_858 ? input_delay_registers_1_13_Re : _GEN_895; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_897 = 5'he == _GEN_858 ? input_delay_registers_1_14_Re : _GEN_896; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_898 = 5'hf == _GEN_858 ? input_delay_registers_1_15_Re : _GEN_897; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_899 = 5'h10 == _GEN_858 ? input_delay_registers_1_16_Re : _GEN_898; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_900 = 5'h11 == _GEN_858 ? input_delay_registers_1_17_Re : _GEN_899; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_901 = 5'h12 == _GEN_858 ? input_delay_registers_1_18_Re : _GEN_900; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_902 = 5'h13 == _GEN_858 ? input_delay_registers_1_19_Re : _GEN_901; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_903 = 5'h14 == _GEN_858 ? input_delay_registers_1_20_Re : _GEN_902; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_904 = 5'h15 == _GEN_858 ? input_delay_registers_1_21_Re : _GEN_903; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_905 = 5'h16 == _GEN_858 ? input_delay_registers_1_22_Re : _GEN_904; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_906 = 5'h17 == _GEN_858 ? input_delay_registers_1_23_Re : _GEN_905; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_916 = 2'h1 == cnt ? 5'h0 : 5'h17; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_917 = 2'h2 == cnt ? 5'h17 : _GEN_916; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_918 = 2'h3 == cnt ? 5'h0 : _GEN_917; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_920 = 5'h1 == _GEN_918 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_921 = 5'h2 == _GEN_918 ? input_delay_registers_1_2_Im : _GEN_920; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_922 = 5'h3 == _GEN_918 ? input_delay_registers_1_3_Im : _GEN_921; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_923 = 5'h4 == _GEN_918 ? input_delay_registers_1_4_Im : _GEN_922; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_924 = 5'h5 == _GEN_918 ? input_delay_registers_1_5_Im : _GEN_923; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_925 = 5'h6 == _GEN_918 ? input_delay_registers_1_6_Im : _GEN_924; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_926 = 5'h7 == _GEN_918 ? input_delay_registers_1_7_Im : _GEN_925; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_927 = 5'h8 == _GEN_918 ? input_delay_registers_1_8_Im : _GEN_926; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_928 = 5'h9 == _GEN_918 ? input_delay_registers_1_9_Im : _GEN_927; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_929 = 5'ha == _GEN_918 ? input_delay_registers_1_10_Im : _GEN_928; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_930 = 5'hb == _GEN_918 ? input_delay_registers_1_11_Im : _GEN_929; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_931 = 5'hc == _GEN_918 ? input_delay_registers_1_12_Im : _GEN_930; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_932 = 5'hd == _GEN_918 ? input_delay_registers_1_13_Im : _GEN_931; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_933 = 5'he == _GEN_918 ? input_delay_registers_1_14_Im : _GEN_932; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_934 = 5'hf == _GEN_918 ? input_delay_registers_1_15_Im : _GEN_933; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_935 = 5'h10 == _GEN_918 ? input_delay_registers_1_16_Im : _GEN_934; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_936 = 5'h11 == _GEN_918 ? input_delay_registers_1_17_Im : _GEN_935; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_937 = 5'h12 == _GEN_918 ? input_delay_registers_1_18_Im : _GEN_936; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_938 = 5'h13 == _GEN_918 ? input_delay_registers_1_19_Im : _GEN_937; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_939 = 5'h14 == _GEN_918 ? input_delay_registers_1_20_Im : _GEN_938; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_940 = 5'h15 == _GEN_918 ? input_delay_registers_1_21_Im : _GEN_939; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_941 = 5'h16 == _GEN_918 ? input_delay_registers_1_22_Im : _GEN_940; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_942 = 5'h17 == _GEN_918 ? input_delay_registers_1_23_Im : _GEN_941; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_944 = 5'h1 == _GEN_918 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_945 = 5'h2 == _GEN_918 ? input_delay_registers_1_2_Re : _GEN_944; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_946 = 5'h3 == _GEN_918 ? input_delay_registers_1_3_Re : _GEN_945; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_947 = 5'h4 == _GEN_918 ? input_delay_registers_1_4_Re : _GEN_946; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_948 = 5'h5 == _GEN_918 ? input_delay_registers_1_5_Re : _GEN_947; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_949 = 5'h6 == _GEN_918 ? input_delay_registers_1_6_Re : _GEN_948; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_950 = 5'h7 == _GEN_918 ? input_delay_registers_1_7_Re : _GEN_949; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_951 = 5'h8 == _GEN_918 ? input_delay_registers_1_8_Re : _GEN_950; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_952 = 5'h9 == _GEN_918 ? input_delay_registers_1_9_Re : _GEN_951; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_953 = 5'ha == _GEN_918 ? input_delay_registers_1_10_Re : _GEN_952; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_954 = 5'hb == _GEN_918 ? input_delay_registers_1_11_Re : _GEN_953; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_955 = 5'hc == _GEN_918 ? input_delay_registers_1_12_Re : _GEN_954; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_956 = 5'hd == _GEN_918 ? input_delay_registers_1_13_Re : _GEN_955; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_957 = 5'he == _GEN_918 ? input_delay_registers_1_14_Re : _GEN_956; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_958 = 5'hf == _GEN_918 ? input_delay_registers_1_15_Re : _GEN_957; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_959 = 5'h10 == _GEN_918 ? input_delay_registers_1_16_Re : _GEN_958; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_960 = 5'h11 == _GEN_918 ? input_delay_registers_1_17_Re : _GEN_959; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_961 = 5'h12 == _GEN_918 ? input_delay_registers_1_18_Re : _GEN_960; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_962 = 5'h13 == _GEN_918 ? input_delay_registers_1_19_Re : _GEN_961; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_963 = 5'h14 == _GEN_918 ? input_delay_registers_1_20_Re : _GEN_962; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_964 = 5'h15 == _GEN_918 ? input_delay_registers_1_21_Re : _GEN_963; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_965 = 5'h16 == _GEN_918 ? input_delay_registers_1_22_Re : _GEN_964; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_966 = 5'h17 == _GEN_918 ? input_delay_registers_1_23_Re : _GEN_965; // @[FFTDesigns.scala 2979:{32,32}]
  wire [2:0] _GEN_972 = 2'h1 == cnt ? 3'h1 : 3'h0; // @[FFTDesigns.scala 2978:{55,55}]
  wire [2:0] _GEN_973 = 2'h2 == cnt ? 3'h3 : _GEN_972; // @[FFTDesigns.scala 2978:{55,55}]
  wire [2:0] _GEN_974 = 2'h3 == cnt ? 3'h4 : _GEN_973; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_2358 = {{1'd0}, _GEN_974}; // @[FFTDesigns.scala 2978:55]
  wire [3:0] _M0_8_in_waddr_0_T_2 = _GEN_2358 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2978:55]
  wire [4:0] _GEN_976 = 2'h1 == cnt ? 5'h0 : 5'h8; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_977 = 2'h2 == cnt ? 5'h8 : _GEN_976; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_978 = 2'h3 == cnt ? 5'h0 : _GEN_977; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_980 = 5'h1 == _GEN_978 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_981 = 5'h2 == _GEN_978 ? input_delay_registers_1_2_Im : _GEN_980; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_982 = 5'h3 == _GEN_978 ? input_delay_registers_1_3_Im : _GEN_981; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_983 = 5'h4 == _GEN_978 ? input_delay_registers_1_4_Im : _GEN_982; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_984 = 5'h5 == _GEN_978 ? input_delay_registers_1_5_Im : _GEN_983; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_985 = 5'h6 == _GEN_978 ? input_delay_registers_1_6_Im : _GEN_984; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_986 = 5'h7 == _GEN_978 ? input_delay_registers_1_7_Im : _GEN_985; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_987 = 5'h8 == _GEN_978 ? input_delay_registers_1_8_Im : _GEN_986; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_988 = 5'h9 == _GEN_978 ? input_delay_registers_1_9_Im : _GEN_987; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_989 = 5'ha == _GEN_978 ? input_delay_registers_1_10_Im : _GEN_988; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_990 = 5'hb == _GEN_978 ? input_delay_registers_1_11_Im : _GEN_989; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_991 = 5'hc == _GEN_978 ? input_delay_registers_1_12_Im : _GEN_990; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_992 = 5'hd == _GEN_978 ? input_delay_registers_1_13_Im : _GEN_991; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_993 = 5'he == _GEN_978 ? input_delay_registers_1_14_Im : _GEN_992; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_994 = 5'hf == _GEN_978 ? input_delay_registers_1_15_Im : _GEN_993; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_995 = 5'h10 == _GEN_978 ? input_delay_registers_1_16_Im : _GEN_994; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_996 = 5'h11 == _GEN_978 ? input_delay_registers_1_17_Im : _GEN_995; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_997 = 5'h12 == _GEN_978 ? input_delay_registers_1_18_Im : _GEN_996; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_998 = 5'h13 == _GEN_978 ? input_delay_registers_1_19_Im : _GEN_997; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_999 = 5'h14 == _GEN_978 ? input_delay_registers_1_20_Im : _GEN_998; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1000 = 5'h15 == _GEN_978 ? input_delay_registers_1_21_Im : _GEN_999; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1001 = 5'h16 == _GEN_978 ? input_delay_registers_1_22_Im : _GEN_1000; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1002 = 5'h17 == _GEN_978 ? input_delay_registers_1_23_Im : _GEN_1001; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1004 = 5'h1 == _GEN_978 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1005 = 5'h2 == _GEN_978 ? input_delay_registers_1_2_Re : _GEN_1004; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1006 = 5'h3 == _GEN_978 ? input_delay_registers_1_3_Re : _GEN_1005; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1007 = 5'h4 == _GEN_978 ? input_delay_registers_1_4_Re : _GEN_1006; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1008 = 5'h5 == _GEN_978 ? input_delay_registers_1_5_Re : _GEN_1007; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1009 = 5'h6 == _GEN_978 ? input_delay_registers_1_6_Re : _GEN_1008; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1010 = 5'h7 == _GEN_978 ? input_delay_registers_1_7_Re : _GEN_1009; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1011 = 5'h8 == _GEN_978 ? input_delay_registers_1_8_Re : _GEN_1010; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1012 = 5'h9 == _GEN_978 ? input_delay_registers_1_9_Re : _GEN_1011; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1013 = 5'ha == _GEN_978 ? input_delay_registers_1_10_Re : _GEN_1012; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1014 = 5'hb == _GEN_978 ? input_delay_registers_1_11_Re : _GEN_1013; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1015 = 5'hc == _GEN_978 ? input_delay_registers_1_12_Re : _GEN_1014; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1016 = 5'hd == _GEN_978 ? input_delay_registers_1_13_Re : _GEN_1015; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1017 = 5'he == _GEN_978 ? input_delay_registers_1_14_Re : _GEN_1016; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1018 = 5'hf == _GEN_978 ? input_delay_registers_1_15_Re : _GEN_1017; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1019 = 5'h10 == _GEN_978 ? input_delay_registers_1_16_Re : _GEN_1018; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1020 = 5'h11 == _GEN_978 ? input_delay_registers_1_17_Re : _GEN_1019; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1021 = 5'h12 == _GEN_978 ? input_delay_registers_1_18_Re : _GEN_1020; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1022 = 5'h13 == _GEN_978 ? input_delay_registers_1_19_Re : _GEN_1021; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1023 = 5'h14 == _GEN_978 ? input_delay_registers_1_20_Re : _GEN_1022; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1024 = 5'h15 == _GEN_978 ? input_delay_registers_1_21_Re : _GEN_1023; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1025 = 5'h16 == _GEN_978 ? input_delay_registers_1_22_Re : _GEN_1024; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1026 = 5'h17 == _GEN_978 ? input_delay_registers_1_23_Re : _GEN_1025; // @[FFTDesigns.scala 2979:{32,32}]
  wire  _GEN_1029 = 2'h2 == cnt ? 1'h0 : 2'h1 == cnt; // @[FFTDesigns.scala 2977:{27,27}]
  wire [2:0] _GEN_1033 = 2'h2 == cnt ? 3'h0 : _GEN_12; // @[FFTDesigns.scala 2978:{55,55}]
  wire [2:0] _GEN_1034 = 2'h3 == cnt ? 3'h5 : _GEN_1033; // @[FFTDesigns.scala 2978:{55,55}]
  wire [3:0] _GEN_2360 = {{1'd0}, _GEN_1034}; // @[FFTDesigns.scala 2978:55]
  wire [3:0] _M0_8_in_waddr_1_T_2 = _GEN_2360 + _M1_0_in_waddr_T; // @[FFTDesigns.scala 2978:55]
  wire [4:0] _GEN_1036 = 2'h1 == cnt ? 5'h10 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1037 = 2'h2 == cnt ? 5'h0 : _GEN_1036; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1038 = 2'h3 == cnt ? 5'h10 : _GEN_1037; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1040 = 5'h1 == _GEN_1038 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1041 = 5'h2 == _GEN_1038 ? input_delay_registers_1_2_Im : _GEN_1040; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1042 = 5'h3 == _GEN_1038 ? input_delay_registers_1_3_Im : _GEN_1041; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1043 = 5'h4 == _GEN_1038 ? input_delay_registers_1_4_Im : _GEN_1042; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1044 = 5'h5 == _GEN_1038 ? input_delay_registers_1_5_Im : _GEN_1043; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1045 = 5'h6 == _GEN_1038 ? input_delay_registers_1_6_Im : _GEN_1044; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1046 = 5'h7 == _GEN_1038 ? input_delay_registers_1_7_Im : _GEN_1045; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1047 = 5'h8 == _GEN_1038 ? input_delay_registers_1_8_Im : _GEN_1046; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1048 = 5'h9 == _GEN_1038 ? input_delay_registers_1_9_Im : _GEN_1047; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1049 = 5'ha == _GEN_1038 ? input_delay_registers_1_10_Im : _GEN_1048; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1050 = 5'hb == _GEN_1038 ? input_delay_registers_1_11_Im : _GEN_1049; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1051 = 5'hc == _GEN_1038 ? input_delay_registers_1_12_Im : _GEN_1050; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1052 = 5'hd == _GEN_1038 ? input_delay_registers_1_13_Im : _GEN_1051; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1053 = 5'he == _GEN_1038 ? input_delay_registers_1_14_Im : _GEN_1052; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1054 = 5'hf == _GEN_1038 ? input_delay_registers_1_15_Im : _GEN_1053; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1055 = 5'h10 == _GEN_1038 ? input_delay_registers_1_16_Im : _GEN_1054; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1056 = 5'h11 == _GEN_1038 ? input_delay_registers_1_17_Im : _GEN_1055; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1057 = 5'h12 == _GEN_1038 ? input_delay_registers_1_18_Im : _GEN_1056; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1058 = 5'h13 == _GEN_1038 ? input_delay_registers_1_19_Im : _GEN_1057; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1059 = 5'h14 == _GEN_1038 ? input_delay_registers_1_20_Im : _GEN_1058; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1060 = 5'h15 == _GEN_1038 ? input_delay_registers_1_21_Im : _GEN_1059; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1061 = 5'h16 == _GEN_1038 ? input_delay_registers_1_22_Im : _GEN_1060; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1062 = 5'h17 == _GEN_1038 ? input_delay_registers_1_23_Im : _GEN_1061; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1064 = 5'h1 == _GEN_1038 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1065 = 5'h2 == _GEN_1038 ? input_delay_registers_1_2_Re : _GEN_1064; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1066 = 5'h3 == _GEN_1038 ? input_delay_registers_1_3_Re : _GEN_1065; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1067 = 5'h4 == _GEN_1038 ? input_delay_registers_1_4_Re : _GEN_1066; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1068 = 5'h5 == _GEN_1038 ? input_delay_registers_1_5_Re : _GEN_1067; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1069 = 5'h6 == _GEN_1038 ? input_delay_registers_1_6_Re : _GEN_1068; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1070 = 5'h7 == _GEN_1038 ? input_delay_registers_1_7_Re : _GEN_1069; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1071 = 5'h8 == _GEN_1038 ? input_delay_registers_1_8_Re : _GEN_1070; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1072 = 5'h9 == _GEN_1038 ? input_delay_registers_1_9_Re : _GEN_1071; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1073 = 5'ha == _GEN_1038 ? input_delay_registers_1_10_Re : _GEN_1072; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1074 = 5'hb == _GEN_1038 ? input_delay_registers_1_11_Re : _GEN_1073; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1075 = 5'hc == _GEN_1038 ? input_delay_registers_1_12_Re : _GEN_1074; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1076 = 5'hd == _GEN_1038 ? input_delay_registers_1_13_Re : _GEN_1075; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1077 = 5'he == _GEN_1038 ? input_delay_registers_1_14_Re : _GEN_1076; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1078 = 5'hf == _GEN_1038 ? input_delay_registers_1_15_Re : _GEN_1077; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1079 = 5'h10 == _GEN_1038 ? input_delay_registers_1_16_Re : _GEN_1078; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1080 = 5'h11 == _GEN_1038 ? input_delay_registers_1_17_Re : _GEN_1079; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1081 = 5'h12 == _GEN_1038 ? input_delay_registers_1_18_Re : _GEN_1080; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1082 = 5'h13 == _GEN_1038 ? input_delay_registers_1_19_Re : _GEN_1081; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1083 = 5'h14 == _GEN_1038 ? input_delay_registers_1_20_Re : _GEN_1082; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1084 = 5'h15 == _GEN_1038 ? input_delay_registers_1_21_Re : _GEN_1083; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1085 = 5'h16 == _GEN_1038 ? input_delay_registers_1_22_Re : _GEN_1084; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1086 = 5'h17 == _GEN_1038 ? input_delay_registers_1_23_Re : _GEN_1085; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1096 = 2'h1 == cnt ? 5'h1 : 5'h9; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1097 = 2'h2 == cnt ? 5'h9 : _GEN_1096; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1098 = 2'h3 == cnt ? 5'h1 : _GEN_1097; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1100 = 5'h1 == _GEN_1098 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1101 = 5'h2 == _GEN_1098 ? input_delay_registers_1_2_Im : _GEN_1100; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1102 = 5'h3 == _GEN_1098 ? input_delay_registers_1_3_Im : _GEN_1101; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1103 = 5'h4 == _GEN_1098 ? input_delay_registers_1_4_Im : _GEN_1102; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1104 = 5'h5 == _GEN_1098 ? input_delay_registers_1_5_Im : _GEN_1103; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1105 = 5'h6 == _GEN_1098 ? input_delay_registers_1_6_Im : _GEN_1104; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1106 = 5'h7 == _GEN_1098 ? input_delay_registers_1_7_Im : _GEN_1105; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1107 = 5'h8 == _GEN_1098 ? input_delay_registers_1_8_Im : _GEN_1106; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1108 = 5'h9 == _GEN_1098 ? input_delay_registers_1_9_Im : _GEN_1107; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1109 = 5'ha == _GEN_1098 ? input_delay_registers_1_10_Im : _GEN_1108; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1110 = 5'hb == _GEN_1098 ? input_delay_registers_1_11_Im : _GEN_1109; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1111 = 5'hc == _GEN_1098 ? input_delay_registers_1_12_Im : _GEN_1110; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1112 = 5'hd == _GEN_1098 ? input_delay_registers_1_13_Im : _GEN_1111; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1113 = 5'he == _GEN_1098 ? input_delay_registers_1_14_Im : _GEN_1112; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1114 = 5'hf == _GEN_1098 ? input_delay_registers_1_15_Im : _GEN_1113; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1115 = 5'h10 == _GEN_1098 ? input_delay_registers_1_16_Im : _GEN_1114; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1116 = 5'h11 == _GEN_1098 ? input_delay_registers_1_17_Im : _GEN_1115; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1117 = 5'h12 == _GEN_1098 ? input_delay_registers_1_18_Im : _GEN_1116; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1118 = 5'h13 == _GEN_1098 ? input_delay_registers_1_19_Im : _GEN_1117; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1119 = 5'h14 == _GEN_1098 ? input_delay_registers_1_20_Im : _GEN_1118; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1120 = 5'h15 == _GEN_1098 ? input_delay_registers_1_21_Im : _GEN_1119; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1121 = 5'h16 == _GEN_1098 ? input_delay_registers_1_22_Im : _GEN_1120; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1122 = 5'h17 == _GEN_1098 ? input_delay_registers_1_23_Im : _GEN_1121; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1124 = 5'h1 == _GEN_1098 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1125 = 5'h2 == _GEN_1098 ? input_delay_registers_1_2_Re : _GEN_1124; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1126 = 5'h3 == _GEN_1098 ? input_delay_registers_1_3_Re : _GEN_1125; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1127 = 5'h4 == _GEN_1098 ? input_delay_registers_1_4_Re : _GEN_1126; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1128 = 5'h5 == _GEN_1098 ? input_delay_registers_1_5_Re : _GEN_1127; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1129 = 5'h6 == _GEN_1098 ? input_delay_registers_1_6_Re : _GEN_1128; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1130 = 5'h7 == _GEN_1098 ? input_delay_registers_1_7_Re : _GEN_1129; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1131 = 5'h8 == _GEN_1098 ? input_delay_registers_1_8_Re : _GEN_1130; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1132 = 5'h9 == _GEN_1098 ? input_delay_registers_1_9_Re : _GEN_1131; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1133 = 5'ha == _GEN_1098 ? input_delay_registers_1_10_Re : _GEN_1132; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1134 = 5'hb == _GEN_1098 ? input_delay_registers_1_11_Re : _GEN_1133; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1135 = 5'hc == _GEN_1098 ? input_delay_registers_1_12_Re : _GEN_1134; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1136 = 5'hd == _GEN_1098 ? input_delay_registers_1_13_Re : _GEN_1135; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1137 = 5'he == _GEN_1098 ? input_delay_registers_1_14_Re : _GEN_1136; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1138 = 5'hf == _GEN_1098 ? input_delay_registers_1_15_Re : _GEN_1137; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1139 = 5'h10 == _GEN_1098 ? input_delay_registers_1_16_Re : _GEN_1138; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1140 = 5'h11 == _GEN_1098 ? input_delay_registers_1_17_Re : _GEN_1139; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1141 = 5'h12 == _GEN_1098 ? input_delay_registers_1_18_Re : _GEN_1140; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1142 = 5'h13 == _GEN_1098 ? input_delay_registers_1_19_Re : _GEN_1141; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1143 = 5'h14 == _GEN_1098 ? input_delay_registers_1_20_Re : _GEN_1142; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1144 = 5'h15 == _GEN_1098 ? input_delay_registers_1_21_Re : _GEN_1143; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1145 = 5'h16 == _GEN_1098 ? input_delay_registers_1_22_Re : _GEN_1144; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1146 = 5'h17 == _GEN_1098 ? input_delay_registers_1_23_Re : _GEN_1145; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1156 = 2'h1 == cnt ? 5'h11 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1157 = 2'h2 == cnt ? 5'h0 : _GEN_1156; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1158 = 2'h3 == cnt ? 5'h11 : _GEN_1157; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1160 = 5'h1 == _GEN_1158 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1161 = 5'h2 == _GEN_1158 ? input_delay_registers_1_2_Im : _GEN_1160; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1162 = 5'h3 == _GEN_1158 ? input_delay_registers_1_3_Im : _GEN_1161; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1163 = 5'h4 == _GEN_1158 ? input_delay_registers_1_4_Im : _GEN_1162; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1164 = 5'h5 == _GEN_1158 ? input_delay_registers_1_5_Im : _GEN_1163; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1165 = 5'h6 == _GEN_1158 ? input_delay_registers_1_6_Im : _GEN_1164; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1166 = 5'h7 == _GEN_1158 ? input_delay_registers_1_7_Im : _GEN_1165; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1167 = 5'h8 == _GEN_1158 ? input_delay_registers_1_8_Im : _GEN_1166; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1168 = 5'h9 == _GEN_1158 ? input_delay_registers_1_9_Im : _GEN_1167; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1169 = 5'ha == _GEN_1158 ? input_delay_registers_1_10_Im : _GEN_1168; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1170 = 5'hb == _GEN_1158 ? input_delay_registers_1_11_Im : _GEN_1169; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1171 = 5'hc == _GEN_1158 ? input_delay_registers_1_12_Im : _GEN_1170; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1172 = 5'hd == _GEN_1158 ? input_delay_registers_1_13_Im : _GEN_1171; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1173 = 5'he == _GEN_1158 ? input_delay_registers_1_14_Im : _GEN_1172; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1174 = 5'hf == _GEN_1158 ? input_delay_registers_1_15_Im : _GEN_1173; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1175 = 5'h10 == _GEN_1158 ? input_delay_registers_1_16_Im : _GEN_1174; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1176 = 5'h11 == _GEN_1158 ? input_delay_registers_1_17_Im : _GEN_1175; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1177 = 5'h12 == _GEN_1158 ? input_delay_registers_1_18_Im : _GEN_1176; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1178 = 5'h13 == _GEN_1158 ? input_delay_registers_1_19_Im : _GEN_1177; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1179 = 5'h14 == _GEN_1158 ? input_delay_registers_1_20_Im : _GEN_1178; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1180 = 5'h15 == _GEN_1158 ? input_delay_registers_1_21_Im : _GEN_1179; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1181 = 5'h16 == _GEN_1158 ? input_delay_registers_1_22_Im : _GEN_1180; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1182 = 5'h17 == _GEN_1158 ? input_delay_registers_1_23_Im : _GEN_1181; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1184 = 5'h1 == _GEN_1158 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1185 = 5'h2 == _GEN_1158 ? input_delay_registers_1_2_Re : _GEN_1184; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1186 = 5'h3 == _GEN_1158 ? input_delay_registers_1_3_Re : _GEN_1185; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1187 = 5'h4 == _GEN_1158 ? input_delay_registers_1_4_Re : _GEN_1186; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1188 = 5'h5 == _GEN_1158 ? input_delay_registers_1_5_Re : _GEN_1187; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1189 = 5'h6 == _GEN_1158 ? input_delay_registers_1_6_Re : _GEN_1188; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1190 = 5'h7 == _GEN_1158 ? input_delay_registers_1_7_Re : _GEN_1189; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1191 = 5'h8 == _GEN_1158 ? input_delay_registers_1_8_Re : _GEN_1190; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1192 = 5'h9 == _GEN_1158 ? input_delay_registers_1_9_Re : _GEN_1191; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1193 = 5'ha == _GEN_1158 ? input_delay_registers_1_10_Re : _GEN_1192; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1194 = 5'hb == _GEN_1158 ? input_delay_registers_1_11_Re : _GEN_1193; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1195 = 5'hc == _GEN_1158 ? input_delay_registers_1_12_Re : _GEN_1194; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1196 = 5'hd == _GEN_1158 ? input_delay_registers_1_13_Re : _GEN_1195; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1197 = 5'he == _GEN_1158 ? input_delay_registers_1_14_Re : _GEN_1196; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1198 = 5'hf == _GEN_1158 ? input_delay_registers_1_15_Re : _GEN_1197; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1199 = 5'h10 == _GEN_1158 ? input_delay_registers_1_16_Re : _GEN_1198; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1200 = 5'h11 == _GEN_1158 ? input_delay_registers_1_17_Re : _GEN_1199; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1201 = 5'h12 == _GEN_1158 ? input_delay_registers_1_18_Re : _GEN_1200; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1202 = 5'h13 == _GEN_1158 ? input_delay_registers_1_19_Re : _GEN_1201; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1203 = 5'h14 == _GEN_1158 ? input_delay_registers_1_20_Re : _GEN_1202; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1204 = 5'h15 == _GEN_1158 ? input_delay_registers_1_21_Re : _GEN_1203; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1205 = 5'h16 == _GEN_1158 ? input_delay_registers_1_22_Re : _GEN_1204; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1206 = 5'h17 == _GEN_1158 ? input_delay_registers_1_23_Re : _GEN_1205; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1216 = 2'h1 == cnt ? 5'h2 : 5'ha; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1217 = 2'h2 == cnt ? 5'ha : _GEN_1216; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1218 = 2'h3 == cnt ? 5'h2 : _GEN_1217; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1220 = 5'h1 == _GEN_1218 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1221 = 5'h2 == _GEN_1218 ? input_delay_registers_1_2_Im : _GEN_1220; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1222 = 5'h3 == _GEN_1218 ? input_delay_registers_1_3_Im : _GEN_1221; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1223 = 5'h4 == _GEN_1218 ? input_delay_registers_1_4_Im : _GEN_1222; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1224 = 5'h5 == _GEN_1218 ? input_delay_registers_1_5_Im : _GEN_1223; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1225 = 5'h6 == _GEN_1218 ? input_delay_registers_1_6_Im : _GEN_1224; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1226 = 5'h7 == _GEN_1218 ? input_delay_registers_1_7_Im : _GEN_1225; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1227 = 5'h8 == _GEN_1218 ? input_delay_registers_1_8_Im : _GEN_1226; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1228 = 5'h9 == _GEN_1218 ? input_delay_registers_1_9_Im : _GEN_1227; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1229 = 5'ha == _GEN_1218 ? input_delay_registers_1_10_Im : _GEN_1228; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1230 = 5'hb == _GEN_1218 ? input_delay_registers_1_11_Im : _GEN_1229; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1231 = 5'hc == _GEN_1218 ? input_delay_registers_1_12_Im : _GEN_1230; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1232 = 5'hd == _GEN_1218 ? input_delay_registers_1_13_Im : _GEN_1231; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1233 = 5'he == _GEN_1218 ? input_delay_registers_1_14_Im : _GEN_1232; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1234 = 5'hf == _GEN_1218 ? input_delay_registers_1_15_Im : _GEN_1233; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1235 = 5'h10 == _GEN_1218 ? input_delay_registers_1_16_Im : _GEN_1234; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1236 = 5'h11 == _GEN_1218 ? input_delay_registers_1_17_Im : _GEN_1235; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1237 = 5'h12 == _GEN_1218 ? input_delay_registers_1_18_Im : _GEN_1236; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1238 = 5'h13 == _GEN_1218 ? input_delay_registers_1_19_Im : _GEN_1237; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1239 = 5'h14 == _GEN_1218 ? input_delay_registers_1_20_Im : _GEN_1238; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1240 = 5'h15 == _GEN_1218 ? input_delay_registers_1_21_Im : _GEN_1239; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1241 = 5'h16 == _GEN_1218 ? input_delay_registers_1_22_Im : _GEN_1240; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1242 = 5'h17 == _GEN_1218 ? input_delay_registers_1_23_Im : _GEN_1241; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1244 = 5'h1 == _GEN_1218 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1245 = 5'h2 == _GEN_1218 ? input_delay_registers_1_2_Re : _GEN_1244; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1246 = 5'h3 == _GEN_1218 ? input_delay_registers_1_3_Re : _GEN_1245; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1247 = 5'h4 == _GEN_1218 ? input_delay_registers_1_4_Re : _GEN_1246; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1248 = 5'h5 == _GEN_1218 ? input_delay_registers_1_5_Re : _GEN_1247; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1249 = 5'h6 == _GEN_1218 ? input_delay_registers_1_6_Re : _GEN_1248; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1250 = 5'h7 == _GEN_1218 ? input_delay_registers_1_7_Re : _GEN_1249; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1251 = 5'h8 == _GEN_1218 ? input_delay_registers_1_8_Re : _GEN_1250; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1252 = 5'h9 == _GEN_1218 ? input_delay_registers_1_9_Re : _GEN_1251; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1253 = 5'ha == _GEN_1218 ? input_delay_registers_1_10_Re : _GEN_1252; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1254 = 5'hb == _GEN_1218 ? input_delay_registers_1_11_Re : _GEN_1253; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1255 = 5'hc == _GEN_1218 ? input_delay_registers_1_12_Re : _GEN_1254; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1256 = 5'hd == _GEN_1218 ? input_delay_registers_1_13_Re : _GEN_1255; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1257 = 5'he == _GEN_1218 ? input_delay_registers_1_14_Re : _GEN_1256; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1258 = 5'hf == _GEN_1218 ? input_delay_registers_1_15_Re : _GEN_1257; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1259 = 5'h10 == _GEN_1218 ? input_delay_registers_1_16_Re : _GEN_1258; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1260 = 5'h11 == _GEN_1218 ? input_delay_registers_1_17_Re : _GEN_1259; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1261 = 5'h12 == _GEN_1218 ? input_delay_registers_1_18_Re : _GEN_1260; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1262 = 5'h13 == _GEN_1218 ? input_delay_registers_1_19_Re : _GEN_1261; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1263 = 5'h14 == _GEN_1218 ? input_delay_registers_1_20_Re : _GEN_1262; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1264 = 5'h15 == _GEN_1218 ? input_delay_registers_1_21_Re : _GEN_1263; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1265 = 5'h16 == _GEN_1218 ? input_delay_registers_1_22_Re : _GEN_1264; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1266 = 5'h17 == _GEN_1218 ? input_delay_registers_1_23_Re : _GEN_1265; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1276 = 2'h1 == cnt ? 5'h12 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1277 = 2'h2 == cnt ? 5'h0 : _GEN_1276; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1278 = 2'h3 == cnt ? 5'h12 : _GEN_1277; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1280 = 5'h1 == _GEN_1278 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1281 = 5'h2 == _GEN_1278 ? input_delay_registers_1_2_Im : _GEN_1280; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1282 = 5'h3 == _GEN_1278 ? input_delay_registers_1_3_Im : _GEN_1281; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1283 = 5'h4 == _GEN_1278 ? input_delay_registers_1_4_Im : _GEN_1282; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1284 = 5'h5 == _GEN_1278 ? input_delay_registers_1_5_Im : _GEN_1283; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1285 = 5'h6 == _GEN_1278 ? input_delay_registers_1_6_Im : _GEN_1284; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1286 = 5'h7 == _GEN_1278 ? input_delay_registers_1_7_Im : _GEN_1285; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1287 = 5'h8 == _GEN_1278 ? input_delay_registers_1_8_Im : _GEN_1286; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1288 = 5'h9 == _GEN_1278 ? input_delay_registers_1_9_Im : _GEN_1287; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1289 = 5'ha == _GEN_1278 ? input_delay_registers_1_10_Im : _GEN_1288; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1290 = 5'hb == _GEN_1278 ? input_delay_registers_1_11_Im : _GEN_1289; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1291 = 5'hc == _GEN_1278 ? input_delay_registers_1_12_Im : _GEN_1290; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1292 = 5'hd == _GEN_1278 ? input_delay_registers_1_13_Im : _GEN_1291; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1293 = 5'he == _GEN_1278 ? input_delay_registers_1_14_Im : _GEN_1292; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1294 = 5'hf == _GEN_1278 ? input_delay_registers_1_15_Im : _GEN_1293; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1295 = 5'h10 == _GEN_1278 ? input_delay_registers_1_16_Im : _GEN_1294; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1296 = 5'h11 == _GEN_1278 ? input_delay_registers_1_17_Im : _GEN_1295; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1297 = 5'h12 == _GEN_1278 ? input_delay_registers_1_18_Im : _GEN_1296; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1298 = 5'h13 == _GEN_1278 ? input_delay_registers_1_19_Im : _GEN_1297; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1299 = 5'h14 == _GEN_1278 ? input_delay_registers_1_20_Im : _GEN_1298; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1300 = 5'h15 == _GEN_1278 ? input_delay_registers_1_21_Im : _GEN_1299; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1301 = 5'h16 == _GEN_1278 ? input_delay_registers_1_22_Im : _GEN_1300; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1302 = 5'h17 == _GEN_1278 ? input_delay_registers_1_23_Im : _GEN_1301; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1304 = 5'h1 == _GEN_1278 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1305 = 5'h2 == _GEN_1278 ? input_delay_registers_1_2_Re : _GEN_1304; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1306 = 5'h3 == _GEN_1278 ? input_delay_registers_1_3_Re : _GEN_1305; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1307 = 5'h4 == _GEN_1278 ? input_delay_registers_1_4_Re : _GEN_1306; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1308 = 5'h5 == _GEN_1278 ? input_delay_registers_1_5_Re : _GEN_1307; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1309 = 5'h6 == _GEN_1278 ? input_delay_registers_1_6_Re : _GEN_1308; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1310 = 5'h7 == _GEN_1278 ? input_delay_registers_1_7_Re : _GEN_1309; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1311 = 5'h8 == _GEN_1278 ? input_delay_registers_1_8_Re : _GEN_1310; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1312 = 5'h9 == _GEN_1278 ? input_delay_registers_1_9_Re : _GEN_1311; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1313 = 5'ha == _GEN_1278 ? input_delay_registers_1_10_Re : _GEN_1312; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1314 = 5'hb == _GEN_1278 ? input_delay_registers_1_11_Re : _GEN_1313; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1315 = 5'hc == _GEN_1278 ? input_delay_registers_1_12_Re : _GEN_1314; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1316 = 5'hd == _GEN_1278 ? input_delay_registers_1_13_Re : _GEN_1315; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1317 = 5'he == _GEN_1278 ? input_delay_registers_1_14_Re : _GEN_1316; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1318 = 5'hf == _GEN_1278 ? input_delay_registers_1_15_Re : _GEN_1317; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1319 = 5'h10 == _GEN_1278 ? input_delay_registers_1_16_Re : _GEN_1318; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1320 = 5'h11 == _GEN_1278 ? input_delay_registers_1_17_Re : _GEN_1319; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1321 = 5'h12 == _GEN_1278 ? input_delay_registers_1_18_Re : _GEN_1320; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1322 = 5'h13 == _GEN_1278 ? input_delay_registers_1_19_Re : _GEN_1321; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1323 = 5'h14 == _GEN_1278 ? input_delay_registers_1_20_Re : _GEN_1322; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1324 = 5'h15 == _GEN_1278 ? input_delay_registers_1_21_Re : _GEN_1323; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1325 = 5'h16 == _GEN_1278 ? input_delay_registers_1_22_Re : _GEN_1324; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1326 = 5'h17 == _GEN_1278 ? input_delay_registers_1_23_Re : _GEN_1325; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1336 = 2'h1 == cnt ? 5'h3 : 5'hb; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1337 = 2'h2 == cnt ? 5'hb : _GEN_1336; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1338 = 2'h3 == cnt ? 5'h3 : _GEN_1337; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1340 = 5'h1 == _GEN_1338 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1341 = 5'h2 == _GEN_1338 ? input_delay_registers_1_2_Im : _GEN_1340; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1342 = 5'h3 == _GEN_1338 ? input_delay_registers_1_3_Im : _GEN_1341; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1343 = 5'h4 == _GEN_1338 ? input_delay_registers_1_4_Im : _GEN_1342; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1344 = 5'h5 == _GEN_1338 ? input_delay_registers_1_5_Im : _GEN_1343; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1345 = 5'h6 == _GEN_1338 ? input_delay_registers_1_6_Im : _GEN_1344; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1346 = 5'h7 == _GEN_1338 ? input_delay_registers_1_7_Im : _GEN_1345; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1347 = 5'h8 == _GEN_1338 ? input_delay_registers_1_8_Im : _GEN_1346; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1348 = 5'h9 == _GEN_1338 ? input_delay_registers_1_9_Im : _GEN_1347; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1349 = 5'ha == _GEN_1338 ? input_delay_registers_1_10_Im : _GEN_1348; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1350 = 5'hb == _GEN_1338 ? input_delay_registers_1_11_Im : _GEN_1349; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1351 = 5'hc == _GEN_1338 ? input_delay_registers_1_12_Im : _GEN_1350; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1352 = 5'hd == _GEN_1338 ? input_delay_registers_1_13_Im : _GEN_1351; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1353 = 5'he == _GEN_1338 ? input_delay_registers_1_14_Im : _GEN_1352; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1354 = 5'hf == _GEN_1338 ? input_delay_registers_1_15_Im : _GEN_1353; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1355 = 5'h10 == _GEN_1338 ? input_delay_registers_1_16_Im : _GEN_1354; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1356 = 5'h11 == _GEN_1338 ? input_delay_registers_1_17_Im : _GEN_1355; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1357 = 5'h12 == _GEN_1338 ? input_delay_registers_1_18_Im : _GEN_1356; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1358 = 5'h13 == _GEN_1338 ? input_delay_registers_1_19_Im : _GEN_1357; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1359 = 5'h14 == _GEN_1338 ? input_delay_registers_1_20_Im : _GEN_1358; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1360 = 5'h15 == _GEN_1338 ? input_delay_registers_1_21_Im : _GEN_1359; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1361 = 5'h16 == _GEN_1338 ? input_delay_registers_1_22_Im : _GEN_1360; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1362 = 5'h17 == _GEN_1338 ? input_delay_registers_1_23_Im : _GEN_1361; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1364 = 5'h1 == _GEN_1338 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1365 = 5'h2 == _GEN_1338 ? input_delay_registers_1_2_Re : _GEN_1364; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1366 = 5'h3 == _GEN_1338 ? input_delay_registers_1_3_Re : _GEN_1365; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1367 = 5'h4 == _GEN_1338 ? input_delay_registers_1_4_Re : _GEN_1366; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1368 = 5'h5 == _GEN_1338 ? input_delay_registers_1_5_Re : _GEN_1367; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1369 = 5'h6 == _GEN_1338 ? input_delay_registers_1_6_Re : _GEN_1368; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1370 = 5'h7 == _GEN_1338 ? input_delay_registers_1_7_Re : _GEN_1369; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1371 = 5'h8 == _GEN_1338 ? input_delay_registers_1_8_Re : _GEN_1370; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1372 = 5'h9 == _GEN_1338 ? input_delay_registers_1_9_Re : _GEN_1371; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1373 = 5'ha == _GEN_1338 ? input_delay_registers_1_10_Re : _GEN_1372; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1374 = 5'hb == _GEN_1338 ? input_delay_registers_1_11_Re : _GEN_1373; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1375 = 5'hc == _GEN_1338 ? input_delay_registers_1_12_Re : _GEN_1374; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1376 = 5'hd == _GEN_1338 ? input_delay_registers_1_13_Re : _GEN_1375; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1377 = 5'he == _GEN_1338 ? input_delay_registers_1_14_Re : _GEN_1376; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1378 = 5'hf == _GEN_1338 ? input_delay_registers_1_15_Re : _GEN_1377; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1379 = 5'h10 == _GEN_1338 ? input_delay_registers_1_16_Re : _GEN_1378; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1380 = 5'h11 == _GEN_1338 ? input_delay_registers_1_17_Re : _GEN_1379; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1381 = 5'h12 == _GEN_1338 ? input_delay_registers_1_18_Re : _GEN_1380; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1382 = 5'h13 == _GEN_1338 ? input_delay_registers_1_19_Re : _GEN_1381; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1383 = 5'h14 == _GEN_1338 ? input_delay_registers_1_20_Re : _GEN_1382; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1384 = 5'h15 == _GEN_1338 ? input_delay_registers_1_21_Re : _GEN_1383; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1385 = 5'h16 == _GEN_1338 ? input_delay_registers_1_22_Re : _GEN_1384; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1386 = 5'h17 == _GEN_1338 ? input_delay_registers_1_23_Re : _GEN_1385; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1396 = 2'h1 == cnt ? 5'h13 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1397 = 2'h2 == cnt ? 5'h0 : _GEN_1396; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1398 = 2'h3 == cnt ? 5'h13 : _GEN_1397; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1400 = 5'h1 == _GEN_1398 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1401 = 5'h2 == _GEN_1398 ? input_delay_registers_1_2_Im : _GEN_1400; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1402 = 5'h3 == _GEN_1398 ? input_delay_registers_1_3_Im : _GEN_1401; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1403 = 5'h4 == _GEN_1398 ? input_delay_registers_1_4_Im : _GEN_1402; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1404 = 5'h5 == _GEN_1398 ? input_delay_registers_1_5_Im : _GEN_1403; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1405 = 5'h6 == _GEN_1398 ? input_delay_registers_1_6_Im : _GEN_1404; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1406 = 5'h7 == _GEN_1398 ? input_delay_registers_1_7_Im : _GEN_1405; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1407 = 5'h8 == _GEN_1398 ? input_delay_registers_1_8_Im : _GEN_1406; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1408 = 5'h9 == _GEN_1398 ? input_delay_registers_1_9_Im : _GEN_1407; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1409 = 5'ha == _GEN_1398 ? input_delay_registers_1_10_Im : _GEN_1408; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1410 = 5'hb == _GEN_1398 ? input_delay_registers_1_11_Im : _GEN_1409; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1411 = 5'hc == _GEN_1398 ? input_delay_registers_1_12_Im : _GEN_1410; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1412 = 5'hd == _GEN_1398 ? input_delay_registers_1_13_Im : _GEN_1411; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1413 = 5'he == _GEN_1398 ? input_delay_registers_1_14_Im : _GEN_1412; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1414 = 5'hf == _GEN_1398 ? input_delay_registers_1_15_Im : _GEN_1413; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1415 = 5'h10 == _GEN_1398 ? input_delay_registers_1_16_Im : _GEN_1414; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1416 = 5'h11 == _GEN_1398 ? input_delay_registers_1_17_Im : _GEN_1415; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1417 = 5'h12 == _GEN_1398 ? input_delay_registers_1_18_Im : _GEN_1416; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1418 = 5'h13 == _GEN_1398 ? input_delay_registers_1_19_Im : _GEN_1417; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1419 = 5'h14 == _GEN_1398 ? input_delay_registers_1_20_Im : _GEN_1418; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1420 = 5'h15 == _GEN_1398 ? input_delay_registers_1_21_Im : _GEN_1419; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1421 = 5'h16 == _GEN_1398 ? input_delay_registers_1_22_Im : _GEN_1420; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1422 = 5'h17 == _GEN_1398 ? input_delay_registers_1_23_Im : _GEN_1421; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1424 = 5'h1 == _GEN_1398 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1425 = 5'h2 == _GEN_1398 ? input_delay_registers_1_2_Re : _GEN_1424; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1426 = 5'h3 == _GEN_1398 ? input_delay_registers_1_3_Re : _GEN_1425; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1427 = 5'h4 == _GEN_1398 ? input_delay_registers_1_4_Re : _GEN_1426; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1428 = 5'h5 == _GEN_1398 ? input_delay_registers_1_5_Re : _GEN_1427; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1429 = 5'h6 == _GEN_1398 ? input_delay_registers_1_6_Re : _GEN_1428; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1430 = 5'h7 == _GEN_1398 ? input_delay_registers_1_7_Re : _GEN_1429; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1431 = 5'h8 == _GEN_1398 ? input_delay_registers_1_8_Re : _GEN_1430; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1432 = 5'h9 == _GEN_1398 ? input_delay_registers_1_9_Re : _GEN_1431; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1433 = 5'ha == _GEN_1398 ? input_delay_registers_1_10_Re : _GEN_1432; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1434 = 5'hb == _GEN_1398 ? input_delay_registers_1_11_Re : _GEN_1433; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1435 = 5'hc == _GEN_1398 ? input_delay_registers_1_12_Re : _GEN_1434; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1436 = 5'hd == _GEN_1398 ? input_delay_registers_1_13_Re : _GEN_1435; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1437 = 5'he == _GEN_1398 ? input_delay_registers_1_14_Re : _GEN_1436; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1438 = 5'hf == _GEN_1398 ? input_delay_registers_1_15_Re : _GEN_1437; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1439 = 5'h10 == _GEN_1398 ? input_delay_registers_1_16_Re : _GEN_1438; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1440 = 5'h11 == _GEN_1398 ? input_delay_registers_1_17_Re : _GEN_1439; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1441 = 5'h12 == _GEN_1398 ? input_delay_registers_1_18_Re : _GEN_1440; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1442 = 5'h13 == _GEN_1398 ? input_delay_registers_1_19_Re : _GEN_1441; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1443 = 5'h14 == _GEN_1398 ? input_delay_registers_1_20_Re : _GEN_1442; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1444 = 5'h15 == _GEN_1398 ? input_delay_registers_1_21_Re : _GEN_1443; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1445 = 5'h16 == _GEN_1398 ? input_delay_registers_1_22_Re : _GEN_1444; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1446 = 5'h17 == _GEN_1398 ? input_delay_registers_1_23_Re : _GEN_1445; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1456 = 2'h1 == cnt ? 5'h4 : 5'hc; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1457 = 2'h2 == cnt ? 5'hc : _GEN_1456; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1458 = 2'h3 == cnt ? 5'h4 : _GEN_1457; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1460 = 5'h1 == _GEN_1458 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1461 = 5'h2 == _GEN_1458 ? input_delay_registers_1_2_Im : _GEN_1460; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1462 = 5'h3 == _GEN_1458 ? input_delay_registers_1_3_Im : _GEN_1461; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1463 = 5'h4 == _GEN_1458 ? input_delay_registers_1_4_Im : _GEN_1462; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1464 = 5'h5 == _GEN_1458 ? input_delay_registers_1_5_Im : _GEN_1463; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1465 = 5'h6 == _GEN_1458 ? input_delay_registers_1_6_Im : _GEN_1464; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1466 = 5'h7 == _GEN_1458 ? input_delay_registers_1_7_Im : _GEN_1465; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1467 = 5'h8 == _GEN_1458 ? input_delay_registers_1_8_Im : _GEN_1466; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1468 = 5'h9 == _GEN_1458 ? input_delay_registers_1_9_Im : _GEN_1467; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1469 = 5'ha == _GEN_1458 ? input_delay_registers_1_10_Im : _GEN_1468; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1470 = 5'hb == _GEN_1458 ? input_delay_registers_1_11_Im : _GEN_1469; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1471 = 5'hc == _GEN_1458 ? input_delay_registers_1_12_Im : _GEN_1470; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1472 = 5'hd == _GEN_1458 ? input_delay_registers_1_13_Im : _GEN_1471; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1473 = 5'he == _GEN_1458 ? input_delay_registers_1_14_Im : _GEN_1472; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1474 = 5'hf == _GEN_1458 ? input_delay_registers_1_15_Im : _GEN_1473; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1475 = 5'h10 == _GEN_1458 ? input_delay_registers_1_16_Im : _GEN_1474; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1476 = 5'h11 == _GEN_1458 ? input_delay_registers_1_17_Im : _GEN_1475; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1477 = 5'h12 == _GEN_1458 ? input_delay_registers_1_18_Im : _GEN_1476; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1478 = 5'h13 == _GEN_1458 ? input_delay_registers_1_19_Im : _GEN_1477; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1479 = 5'h14 == _GEN_1458 ? input_delay_registers_1_20_Im : _GEN_1478; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1480 = 5'h15 == _GEN_1458 ? input_delay_registers_1_21_Im : _GEN_1479; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1481 = 5'h16 == _GEN_1458 ? input_delay_registers_1_22_Im : _GEN_1480; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1482 = 5'h17 == _GEN_1458 ? input_delay_registers_1_23_Im : _GEN_1481; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1484 = 5'h1 == _GEN_1458 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1485 = 5'h2 == _GEN_1458 ? input_delay_registers_1_2_Re : _GEN_1484; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1486 = 5'h3 == _GEN_1458 ? input_delay_registers_1_3_Re : _GEN_1485; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1487 = 5'h4 == _GEN_1458 ? input_delay_registers_1_4_Re : _GEN_1486; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1488 = 5'h5 == _GEN_1458 ? input_delay_registers_1_5_Re : _GEN_1487; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1489 = 5'h6 == _GEN_1458 ? input_delay_registers_1_6_Re : _GEN_1488; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1490 = 5'h7 == _GEN_1458 ? input_delay_registers_1_7_Re : _GEN_1489; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1491 = 5'h8 == _GEN_1458 ? input_delay_registers_1_8_Re : _GEN_1490; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1492 = 5'h9 == _GEN_1458 ? input_delay_registers_1_9_Re : _GEN_1491; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1493 = 5'ha == _GEN_1458 ? input_delay_registers_1_10_Re : _GEN_1492; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1494 = 5'hb == _GEN_1458 ? input_delay_registers_1_11_Re : _GEN_1493; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1495 = 5'hc == _GEN_1458 ? input_delay_registers_1_12_Re : _GEN_1494; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1496 = 5'hd == _GEN_1458 ? input_delay_registers_1_13_Re : _GEN_1495; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1497 = 5'he == _GEN_1458 ? input_delay_registers_1_14_Re : _GEN_1496; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1498 = 5'hf == _GEN_1458 ? input_delay_registers_1_15_Re : _GEN_1497; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1499 = 5'h10 == _GEN_1458 ? input_delay_registers_1_16_Re : _GEN_1498; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1500 = 5'h11 == _GEN_1458 ? input_delay_registers_1_17_Re : _GEN_1499; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1501 = 5'h12 == _GEN_1458 ? input_delay_registers_1_18_Re : _GEN_1500; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1502 = 5'h13 == _GEN_1458 ? input_delay_registers_1_19_Re : _GEN_1501; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1503 = 5'h14 == _GEN_1458 ? input_delay_registers_1_20_Re : _GEN_1502; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1504 = 5'h15 == _GEN_1458 ? input_delay_registers_1_21_Re : _GEN_1503; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1505 = 5'h16 == _GEN_1458 ? input_delay_registers_1_22_Re : _GEN_1504; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1506 = 5'h17 == _GEN_1458 ? input_delay_registers_1_23_Re : _GEN_1505; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1516 = 2'h1 == cnt ? 5'h14 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1517 = 2'h2 == cnt ? 5'h0 : _GEN_1516; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1518 = 2'h3 == cnt ? 5'h14 : _GEN_1517; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1520 = 5'h1 == _GEN_1518 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1521 = 5'h2 == _GEN_1518 ? input_delay_registers_1_2_Im : _GEN_1520; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1522 = 5'h3 == _GEN_1518 ? input_delay_registers_1_3_Im : _GEN_1521; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1523 = 5'h4 == _GEN_1518 ? input_delay_registers_1_4_Im : _GEN_1522; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1524 = 5'h5 == _GEN_1518 ? input_delay_registers_1_5_Im : _GEN_1523; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1525 = 5'h6 == _GEN_1518 ? input_delay_registers_1_6_Im : _GEN_1524; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1526 = 5'h7 == _GEN_1518 ? input_delay_registers_1_7_Im : _GEN_1525; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1527 = 5'h8 == _GEN_1518 ? input_delay_registers_1_8_Im : _GEN_1526; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1528 = 5'h9 == _GEN_1518 ? input_delay_registers_1_9_Im : _GEN_1527; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1529 = 5'ha == _GEN_1518 ? input_delay_registers_1_10_Im : _GEN_1528; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1530 = 5'hb == _GEN_1518 ? input_delay_registers_1_11_Im : _GEN_1529; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1531 = 5'hc == _GEN_1518 ? input_delay_registers_1_12_Im : _GEN_1530; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1532 = 5'hd == _GEN_1518 ? input_delay_registers_1_13_Im : _GEN_1531; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1533 = 5'he == _GEN_1518 ? input_delay_registers_1_14_Im : _GEN_1532; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1534 = 5'hf == _GEN_1518 ? input_delay_registers_1_15_Im : _GEN_1533; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1535 = 5'h10 == _GEN_1518 ? input_delay_registers_1_16_Im : _GEN_1534; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1536 = 5'h11 == _GEN_1518 ? input_delay_registers_1_17_Im : _GEN_1535; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1537 = 5'h12 == _GEN_1518 ? input_delay_registers_1_18_Im : _GEN_1536; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1538 = 5'h13 == _GEN_1518 ? input_delay_registers_1_19_Im : _GEN_1537; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1539 = 5'h14 == _GEN_1518 ? input_delay_registers_1_20_Im : _GEN_1538; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1540 = 5'h15 == _GEN_1518 ? input_delay_registers_1_21_Im : _GEN_1539; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1541 = 5'h16 == _GEN_1518 ? input_delay_registers_1_22_Im : _GEN_1540; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1542 = 5'h17 == _GEN_1518 ? input_delay_registers_1_23_Im : _GEN_1541; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1544 = 5'h1 == _GEN_1518 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1545 = 5'h2 == _GEN_1518 ? input_delay_registers_1_2_Re : _GEN_1544; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1546 = 5'h3 == _GEN_1518 ? input_delay_registers_1_3_Re : _GEN_1545; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1547 = 5'h4 == _GEN_1518 ? input_delay_registers_1_4_Re : _GEN_1546; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1548 = 5'h5 == _GEN_1518 ? input_delay_registers_1_5_Re : _GEN_1547; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1549 = 5'h6 == _GEN_1518 ? input_delay_registers_1_6_Re : _GEN_1548; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1550 = 5'h7 == _GEN_1518 ? input_delay_registers_1_7_Re : _GEN_1549; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1551 = 5'h8 == _GEN_1518 ? input_delay_registers_1_8_Re : _GEN_1550; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1552 = 5'h9 == _GEN_1518 ? input_delay_registers_1_9_Re : _GEN_1551; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1553 = 5'ha == _GEN_1518 ? input_delay_registers_1_10_Re : _GEN_1552; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1554 = 5'hb == _GEN_1518 ? input_delay_registers_1_11_Re : _GEN_1553; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1555 = 5'hc == _GEN_1518 ? input_delay_registers_1_12_Re : _GEN_1554; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1556 = 5'hd == _GEN_1518 ? input_delay_registers_1_13_Re : _GEN_1555; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1557 = 5'he == _GEN_1518 ? input_delay_registers_1_14_Re : _GEN_1556; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1558 = 5'hf == _GEN_1518 ? input_delay_registers_1_15_Re : _GEN_1557; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1559 = 5'h10 == _GEN_1518 ? input_delay_registers_1_16_Re : _GEN_1558; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1560 = 5'h11 == _GEN_1518 ? input_delay_registers_1_17_Re : _GEN_1559; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1561 = 5'h12 == _GEN_1518 ? input_delay_registers_1_18_Re : _GEN_1560; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1562 = 5'h13 == _GEN_1518 ? input_delay_registers_1_19_Re : _GEN_1561; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1563 = 5'h14 == _GEN_1518 ? input_delay_registers_1_20_Re : _GEN_1562; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1564 = 5'h15 == _GEN_1518 ? input_delay_registers_1_21_Re : _GEN_1563; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1565 = 5'h16 == _GEN_1518 ? input_delay_registers_1_22_Re : _GEN_1564; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1566 = 5'h17 == _GEN_1518 ? input_delay_registers_1_23_Re : _GEN_1565; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1576 = 2'h1 == cnt ? 5'h5 : 5'hd; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1577 = 2'h2 == cnt ? 5'hd : _GEN_1576; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1578 = 2'h3 == cnt ? 5'h5 : _GEN_1577; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1580 = 5'h1 == _GEN_1578 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1581 = 5'h2 == _GEN_1578 ? input_delay_registers_1_2_Im : _GEN_1580; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1582 = 5'h3 == _GEN_1578 ? input_delay_registers_1_3_Im : _GEN_1581; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1583 = 5'h4 == _GEN_1578 ? input_delay_registers_1_4_Im : _GEN_1582; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1584 = 5'h5 == _GEN_1578 ? input_delay_registers_1_5_Im : _GEN_1583; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1585 = 5'h6 == _GEN_1578 ? input_delay_registers_1_6_Im : _GEN_1584; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1586 = 5'h7 == _GEN_1578 ? input_delay_registers_1_7_Im : _GEN_1585; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1587 = 5'h8 == _GEN_1578 ? input_delay_registers_1_8_Im : _GEN_1586; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1588 = 5'h9 == _GEN_1578 ? input_delay_registers_1_9_Im : _GEN_1587; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1589 = 5'ha == _GEN_1578 ? input_delay_registers_1_10_Im : _GEN_1588; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1590 = 5'hb == _GEN_1578 ? input_delay_registers_1_11_Im : _GEN_1589; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1591 = 5'hc == _GEN_1578 ? input_delay_registers_1_12_Im : _GEN_1590; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1592 = 5'hd == _GEN_1578 ? input_delay_registers_1_13_Im : _GEN_1591; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1593 = 5'he == _GEN_1578 ? input_delay_registers_1_14_Im : _GEN_1592; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1594 = 5'hf == _GEN_1578 ? input_delay_registers_1_15_Im : _GEN_1593; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1595 = 5'h10 == _GEN_1578 ? input_delay_registers_1_16_Im : _GEN_1594; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1596 = 5'h11 == _GEN_1578 ? input_delay_registers_1_17_Im : _GEN_1595; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1597 = 5'h12 == _GEN_1578 ? input_delay_registers_1_18_Im : _GEN_1596; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1598 = 5'h13 == _GEN_1578 ? input_delay_registers_1_19_Im : _GEN_1597; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1599 = 5'h14 == _GEN_1578 ? input_delay_registers_1_20_Im : _GEN_1598; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1600 = 5'h15 == _GEN_1578 ? input_delay_registers_1_21_Im : _GEN_1599; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1601 = 5'h16 == _GEN_1578 ? input_delay_registers_1_22_Im : _GEN_1600; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1602 = 5'h17 == _GEN_1578 ? input_delay_registers_1_23_Im : _GEN_1601; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1604 = 5'h1 == _GEN_1578 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1605 = 5'h2 == _GEN_1578 ? input_delay_registers_1_2_Re : _GEN_1604; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1606 = 5'h3 == _GEN_1578 ? input_delay_registers_1_3_Re : _GEN_1605; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1607 = 5'h4 == _GEN_1578 ? input_delay_registers_1_4_Re : _GEN_1606; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1608 = 5'h5 == _GEN_1578 ? input_delay_registers_1_5_Re : _GEN_1607; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1609 = 5'h6 == _GEN_1578 ? input_delay_registers_1_6_Re : _GEN_1608; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1610 = 5'h7 == _GEN_1578 ? input_delay_registers_1_7_Re : _GEN_1609; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1611 = 5'h8 == _GEN_1578 ? input_delay_registers_1_8_Re : _GEN_1610; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1612 = 5'h9 == _GEN_1578 ? input_delay_registers_1_9_Re : _GEN_1611; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1613 = 5'ha == _GEN_1578 ? input_delay_registers_1_10_Re : _GEN_1612; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1614 = 5'hb == _GEN_1578 ? input_delay_registers_1_11_Re : _GEN_1613; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1615 = 5'hc == _GEN_1578 ? input_delay_registers_1_12_Re : _GEN_1614; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1616 = 5'hd == _GEN_1578 ? input_delay_registers_1_13_Re : _GEN_1615; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1617 = 5'he == _GEN_1578 ? input_delay_registers_1_14_Re : _GEN_1616; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1618 = 5'hf == _GEN_1578 ? input_delay_registers_1_15_Re : _GEN_1617; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1619 = 5'h10 == _GEN_1578 ? input_delay_registers_1_16_Re : _GEN_1618; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1620 = 5'h11 == _GEN_1578 ? input_delay_registers_1_17_Re : _GEN_1619; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1621 = 5'h12 == _GEN_1578 ? input_delay_registers_1_18_Re : _GEN_1620; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1622 = 5'h13 == _GEN_1578 ? input_delay_registers_1_19_Re : _GEN_1621; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1623 = 5'h14 == _GEN_1578 ? input_delay_registers_1_20_Re : _GEN_1622; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1624 = 5'h15 == _GEN_1578 ? input_delay_registers_1_21_Re : _GEN_1623; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1625 = 5'h16 == _GEN_1578 ? input_delay_registers_1_22_Re : _GEN_1624; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1626 = 5'h17 == _GEN_1578 ? input_delay_registers_1_23_Re : _GEN_1625; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1636 = 2'h1 == cnt ? 5'h15 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1637 = 2'h2 == cnt ? 5'h0 : _GEN_1636; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1638 = 2'h3 == cnt ? 5'h15 : _GEN_1637; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1640 = 5'h1 == _GEN_1638 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1641 = 5'h2 == _GEN_1638 ? input_delay_registers_1_2_Im : _GEN_1640; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1642 = 5'h3 == _GEN_1638 ? input_delay_registers_1_3_Im : _GEN_1641; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1643 = 5'h4 == _GEN_1638 ? input_delay_registers_1_4_Im : _GEN_1642; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1644 = 5'h5 == _GEN_1638 ? input_delay_registers_1_5_Im : _GEN_1643; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1645 = 5'h6 == _GEN_1638 ? input_delay_registers_1_6_Im : _GEN_1644; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1646 = 5'h7 == _GEN_1638 ? input_delay_registers_1_7_Im : _GEN_1645; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1647 = 5'h8 == _GEN_1638 ? input_delay_registers_1_8_Im : _GEN_1646; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1648 = 5'h9 == _GEN_1638 ? input_delay_registers_1_9_Im : _GEN_1647; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1649 = 5'ha == _GEN_1638 ? input_delay_registers_1_10_Im : _GEN_1648; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1650 = 5'hb == _GEN_1638 ? input_delay_registers_1_11_Im : _GEN_1649; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1651 = 5'hc == _GEN_1638 ? input_delay_registers_1_12_Im : _GEN_1650; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1652 = 5'hd == _GEN_1638 ? input_delay_registers_1_13_Im : _GEN_1651; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1653 = 5'he == _GEN_1638 ? input_delay_registers_1_14_Im : _GEN_1652; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1654 = 5'hf == _GEN_1638 ? input_delay_registers_1_15_Im : _GEN_1653; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1655 = 5'h10 == _GEN_1638 ? input_delay_registers_1_16_Im : _GEN_1654; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1656 = 5'h11 == _GEN_1638 ? input_delay_registers_1_17_Im : _GEN_1655; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1657 = 5'h12 == _GEN_1638 ? input_delay_registers_1_18_Im : _GEN_1656; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1658 = 5'h13 == _GEN_1638 ? input_delay_registers_1_19_Im : _GEN_1657; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1659 = 5'h14 == _GEN_1638 ? input_delay_registers_1_20_Im : _GEN_1658; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1660 = 5'h15 == _GEN_1638 ? input_delay_registers_1_21_Im : _GEN_1659; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1661 = 5'h16 == _GEN_1638 ? input_delay_registers_1_22_Im : _GEN_1660; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1662 = 5'h17 == _GEN_1638 ? input_delay_registers_1_23_Im : _GEN_1661; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1664 = 5'h1 == _GEN_1638 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1665 = 5'h2 == _GEN_1638 ? input_delay_registers_1_2_Re : _GEN_1664; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1666 = 5'h3 == _GEN_1638 ? input_delay_registers_1_3_Re : _GEN_1665; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1667 = 5'h4 == _GEN_1638 ? input_delay_registers_1_4_Re : _GEN_1666; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1668 = 5'h5 == _GEN_1638 ? input_delay_registers_1_5_Re : _GEN_1667; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1669 = 5'h6 == _GEN_1638 ? input_delay_registers_1_6_Re : _GEN_1668; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1670 = 5'h7 == _GEN_1638 ? input_delay_registers_1_7_Re : _GEN_1669; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1671 = 5'h8 == _GEN_1638 ? input_delay_registers_1_8_Re : _GEN_1670; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1672 = 5'h9 == _GEN_1638 ? input_delay_registers_1_9_Re : _GEN_1671; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1673 = 5'ha == _GEN_1638 ? input_delay_registers_1_10_Re : _GEN_1672; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1674 = 5'hb == _GEN_1638 ? input_delay_registers_1_11_Re : _GEN_1673; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1675 = 5'hc == _GEN_1638 ? input_delay_registers_1_12_Re : _GEN_1674; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1676 = 5'hd == _GEN_1638 ? input_delay_registers_1_13_Re : _GEN_1675; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1677 = 5'he == _GEN_1638 ? input_delay_registers_1_14_Re : _GEN_1676; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1678 = 5'hf == _GEN_1638 ? input_delay_registers_1_15_Re : _GEN_1677; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1679 = 5'h10 == _GEN_1638 ? input_delay_registers_1_16_Re : _GEN_1678; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1680 = 5'h11 == _GEN_1638 ? input_delay_registers_1_17_Re : _GEN_1679; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1681 = 5'h12 == _GEN_1638 ? input_delay_registers_1_18_Re : _GEN_1680; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1682 = 5'h13 == _GEN_1638 ? input_delay_registers_1_19_Re : _GEN_1681; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1683 = 5'h14 == _GEN_1638 ? input_delay_registers_1_20_Re : _GEN_1682; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1684 = 5'h15 == _GEN_1638 ? input_delay_registers_1_21_Re : _GEN_1683; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1685 = 5'h16 == _GEN_1638 ? input_delay_registers_1_22_Re : _GEN_1684; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1686 = 5'h17 == _GEN_1638 ? input_delay_registers_1_23_Re : _GEN_1685; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1696 = 2'h1 == cnt ? 5'h6 : 5'he; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1697 = 2'h2 == cnt ? 5'he : _GEN_1696; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1698 = 2'h3 == cnt ? 5'h6 : _GEN_1697; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1700 = 5'h1 == _GEN_1698 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1701 = 5'h2 == _GEN_1698 ? input_delay_registers_1_2_Im : _GEN_1700; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1702 = 5'h3 == _GEN_1698 ? input_delay_registers_1_3_Im : _GEN_1701; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1703 = 5'h4 == _GEN_1698 ? input_delay_registers_1_4_Im : _GEN_1702; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1704 = 5'h5 == _GEN_1698 ? input_delay_registers_1_5_Im : _GEN_1703; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1705 = 5'h6 == _GEN_1698 ? input_delay_registers_1_6_Im : _GEN_1704; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1706 = 5'h7 == _GEN_1698 ? input_delay_registers_1_7_Im : _GEN_1705; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1707 = 5'h8 == _GEN_1698 ? input_delay_registers_1_8_Im : _GEN_1706; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1708 = 5'h9 == _GEN_1698 ? input_delay_registers_1_9_Im : _GEN_1707; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1709 = 5'ha == _GEN_1698 ? input_delay_registers_1_10_Im : _GEN_1708; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1710 = 5'hb == _GEN_1698 ? input_delay_registers_1_11_Im : _GEN_1709; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1711 = 5'hc == _GEN_1698 ? input_delay_registers_1_12_Im : _GEN_1710; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1712 = 5'hd == _GEN_1698 ? input_delay_registers_1_13_Im : _GEN_1711; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1713 = 5'he == _GEN_1698 ? input_delay_registers_1_14_Im : _GEN_1712; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1714 = 5'hf == _GEN_1698 ? input_delay_registers_1_15_Im : _GEN_1713; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1715 = 5'h10 == _GEN_1698 ? input_delay_registers_1_16_Im : _GEN_1714; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1716 = 5'h11 == _GEN_1698 ? input_delay_registers_1_17_Im : _GEN_1715; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1717 = 5'h12 == _GEN_1698 ? input_delay_registers_1_18_Im : _GEN_1716; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1718 = 5'h13 == _GEN_1698 ? input_delay_registers_1_19_Im : _GEN_1717; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1719 = 5'h14 == _GEN_1698 ? input_delay_registers_1_20_Im : _GEN_1718; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1720 = 5'h15 == _GEN_1698 ? input_delay_registers_1_21_Im : _GEN_1719; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1721 = 5'h16 == _GEN_1698 ? input_delay_registers_1_22_Im : _GEN_1720; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1722 = 5'h17 == _GEN_1698 ? input_delay_registers_1_23_Im : _GEN_1721; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1724 = 5'h1 == _GEN_1698 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1725 = 5'h2 == _GEN_1698 ? input_delay_registers_1_2_Re : _GEN_1724; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1726 = 5'h3 == _GEN_1698 ? input_delay_registers_1_3_Re : _GEN_1725; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1727 = 5'h4 == _GEN_1698 ? input_delay_registers_1_4_Re : _GEN_1726; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1728 = 5'h5 == _GEN_1698 ? input_delay_registers_1_5_Re : _GEN_1727; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1729 = 5'h6 == _GEN_1698 ? input_delay_registers_1_6_Re : _GEN_1728; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1730 = 5'h7 == _GEN_1698 ? input_delay_registers_1_7_Re : _GEN_1729; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1731 = 5'h8 == _GEN_1698 ? input_delay_registers_1_8_Re : _GEN_1730; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1732 = 5'h9 == _GEN_1698 ? input_delay_registers_1_9_Re : _GEN_1731; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1733 = 5'ha == _GEN_1698 ? input_delay_registers_1_10_Re : _GEN_1732; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1734 = 5'hb == _GEN_1698 ? input_delay_registers_1_11_Re : _GEN_1733; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1735 = 5'hc == _GEN_1698 ? input_delay_registers_1_12_Re : _GEN_1734; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1736 = 5'hd == _GEN_1698 ? input_delay_registers_1_13_Re : _GEN_1735; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1737 = 5'he == _GEN_1698 ? input_delay_registers_1_14_Re : _GEN_1736; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1738 = 5'hf == _GEN_1698 ? input_delay_registers_1_15_Re : _GEN_1737; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1739 = 5'h10 == _GEN_1698 ? input_delay_registers_1_16_Re : _GEN_1738; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1740 = 5'h11 == _GEN_1698 ? input_delay_registers_1_17_Re : _GEN_1739; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1741 = 5'h12 == _GEN_1698 ? input_delay_registers_1_18_Re : _GEN_1740; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1742 = 5'h13 == _GEN_1698 ? input_delay_registers_1_19_Re : _GEN_1741; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1743 = 5'h14 == _GEN_1698 ? input_delay_registers_1_20_Re : _GEN_1742; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1744 = 5'h15 == _GEN_1698 ? input_delay_registers_1_21_Re : _GEN_1743; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1745 = 5'h16 == _GEN_1698 ? input_delay_registers_1_22_Re : _GEN_1744; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1746 = 5'h17 == _GEN_1698 ? input_delay_registers_1_23_Re : _GEN_1745; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1756 = 2'h1 == cnt ? 5'h16 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1757 = 2'h2 == cnt ? 5'h0 : _GEN_1756; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1758 = 2'h3 == cnt ? 5'h16 : _GEN_1757; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1760 = 5'h1 == _GEN_1758 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1761 = 5'h2 == _GEN_1758 ? input_delay_registers_1_2_Im : _GEN_1760; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1762 = 5'h3 == _GEN_1758 ? input_delay_registers_1_3_Im : _GEN_1761; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1763 = 5'h4 == _GEN_1758 ? input_delay_registers_1_4_Im : _GEN_1762; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1764 = 5'h5 == _GEN_1758 ? input_delay_registers_1_5_Im : _GEN_1763; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1765 = 5'h6 == _GEN_1758 ? input_delay_registers_1_6_Im : _GEN_1764; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1766 = 5'h7 == _GEN_1758 ? input_delay_registers_1_7_Im : _GEN_1765; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1767 = 5'h8 == _GEN_1758 ? input_delay_registers_1_8_Im : _GEN_1766; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1768 = 5'h9 == _GEN_1758 ? input_delay_registers_1_9_Im : _GEN_1767; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1769 = 5'ha == _GEN_1758 ? input_delay_registers_1_10_Im : _GEN_1768; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1770 = 5'hb == _GEN_1758 ? input_delay_registers_1_11_Im : _GEN_1769; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1771 = 5'hc == _GEN_1758 ? input_delay_registers_1_12_Im : _GEN_1770; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1772 = 5'hd == _GEN_1758 ? input_delay_registers_1_13_Im : _GEN_1771; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1773 = 5'he == _GEN_1758 ? input_delay_registers_1_14_Im : _GEN_1772; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1774 = 5'hf == _GEN_1758 ? input_delay_registers_1_15_Im : _GEN_1773; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1775 = 5'h10 == _GEN_1758 ? input_delay_registers_1_16_Im : _GEN_1774; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1776 = 5'h11 == _GEN_1758 ? input_delay_registers_1_17_Im : _GEN_1775; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1777 = 5'h12 == _GEN_1758 ? input_delay_registers_1_18_Im : _GEN_1776; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1778 = 5'h13 == _GEN_1758 ? input_delay_registers_1_19_Im : _GEN_1777; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1779 = 5'h14 == _GEN_1758 ? input_delay_registers_1_20_Im : _GEN_1778; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1780 = 5'h15 == _GEN_1758 ? input_delay_registers_1_21_Im : _GEN_1779; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1781 = 5'h16 == _GEN_1758 ? input_delay_registers_1_22_Im : _GEN_1780; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1782 = 5'h17 == _GEN_1758 ? input_delay_registers_1_23_Im : _GEN_1781; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1784 = 5'h1 == _GEN_1758 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1785 = 5'h2 == _GEN_1758 ? input_delay_registers_1_2_Re : _GEN_1784; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1786 = 5'h3 == _GEN_1758 ? input_delay_registers_1_3_Re : _GEN_1785; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1787 = 5'h4 == _GEN_1758 ? input_delay_registers_1_4_Re : _GEN_1786; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1788 = 5'h5 == _GEN_1758 ? input_delay_registers_1_5_Re : _GEN_1787; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1789 = 5'h6 == _GEN_1758 ? input_delay_registers_1_6_Re : _GEN_1788; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1790 = 5'h7 == _GEN_1758 ? input_delay_registers_1_7_Re : _GEN_1789; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1791 = 5'h8 == _GEN_1758 ? input_delay_registers_1_8_Re : _GEN_1790; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1792 = 5'h9 == _GEN_1758 ? input_delay_registers_1_9_Re : _GEN_1791; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1793 = 5'ha == _GEN_1758 ? input_delay_registers_1_10_Re : _GEN_1792; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1794 = 5'hb == _GEN_1758 ? input_delay_registers_1_11_Re : _GEN_1793; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1795 = 5'hc == _GEN_1758 ? input_delay_registers_1_12_Re : _GEN_1794; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1796 = 5'hd == _GEN_1758 ? input_delay_registers_1_13_Re : _GEN_1795; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1797 = 5'he == _GEN_1758 ? input_delay_registers_1_14_Re : _GEN_1796; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1798 = 5'hf == _GEN_1758 ? input_delay_registers_1_15_Re : _GEN_1797; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1799 = 5'h10 == _GEN_1758 ? input_delay_registers_1_16_Re : _GEN_1798; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1800 = 5'h11 == _GEN_1758 ? input_delay_registers_1_17_Re : _GEN_1799; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1801 = 5'h12 == _GEN_1758 ? input_delay_registers_1_18_Re : _GEN_1800; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1802 = 5'h13 == _GEN_1758 ? input_delay_registers_1_19_Re : _GEN_1801; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1803 = 5'h14 == _GEN_1758 ? input_delay_registers_1_20_Re : _GEN_1802; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1804 = 5'h15 == _GEN_1758 ? input_delay_registers_1_21_Re : _GEN_1803; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1805 = 5'h16 == _GEN_1758 ? input_delay_registers_1_22_Re : _GEN_1804; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1806 = 5'h17 == _GEN_1758 ? input_delay_registers_1_23_Re : _GEN_1805; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1816 = 2'h1 == cnt ? 5'h7 : 5'hf; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1817 = 2'h2 == cnt ? 5'hf : _GEN_1816; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1818 = 2'h3 == cnt ? 5'h7 : _GEN_1817; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1820 = 5'h1 == _GEN_1818 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1821 = 5'h2 == _GEN_1818 ? input_delay_registers_1_2_Im : _GEN_1820; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1822 = 5'h3 == _GEN_1818 ? input_delay_registers_1_3_Im : _GEN_1821; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1823 = 5'h4 == _GEN_1818 ? input_delay_registers_1_4_Im : _GEN_1822; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1824 = 5'h5 == _GEN_1818 ? input_delay_registers_1_5_Im : _GEN_1823; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1825 = 5'h6 == _GEN_1818 ? input_delay_registers_1_6_Im : _GEN_1824; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1826 = 5'h7 == _GEN_1818 ? input_delay_registers_1_7_Im : _GEN_1825; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1827 = 5'h8 == _GEN_1818 ? input_delay_registers_1_8_Im : _GEN_1826; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1828 = 5'h9 == _GEN_1818 ? input_delay_registers_1_9_Im : _GEN_1827; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1829 = 5'ha == _GEN_1818 ? input_delay_registers_1_10_Im : _GEN_1828; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1830 = 5'hb == _GEN_1818 ? input_delay_registers_1_11_Im : _GEN_1829; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1831 = 5'hc == _GEN_1818 ? input_delay_registers_1_12_Im : _GEN_1830; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1832 = 5'hd == _GEN_1818 ? input_delay_registers_1_13_Im : _GEN_1831; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1833 = 5'he == _GEN_1818 ? input_delay_registers_1_14_Im : _GEN_1832; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1834 = 5'hf == _GEN_1818 ? input_delay_registers_1_15_Im : _GEN_1833; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1835 = 5'h10 == _GEN_1818 ? input_delay_registers_1_16_Im : _GEN_1834; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1836 = 5'h11 == _GEN_1818 ? input_delay_registers_1_17_Im : _GEN_1835; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1837 = 5'h12 == _GEN_1818 ? input_delay_registers_1_18_Im : _GEN_1836; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1838 = 5'h13 == _GEN_1818 ? input_delay_registers_1_19_Im : _GEN_1837; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1839 = 5'h14 == _GEN_1818 ? input_delay_registers_1_20_Im : _GEN_1838; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1840 = 5'h15 == _GEN_1818 ? input_delay_registers_1_21_Im : _GEN_1839; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1841 = 5'h16 == _GEN_1818 ? input_delay_registers_1_22_Im : _GEN_1840; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1842 = 5'h17 == _GEN_1818 ? input_delay_registers_1_23_Im : _GEN_1841; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1844 = 5'h1 == _GEN_1818 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1845 = 5'h2 == _GEN_1818 ? input_delay_registers_1_2_Re : _GEN_1844; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1846 = 5'h3 == _GEN_1818 ? input_delay_registers_1_3_Re : _GEN_1845; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1847 = 5'h4 == _GEN_1818 ? input_delay_registers_1_4_Re : _GEN_1846; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1848 = 5'h5 == _GEN_1818 ? input_delay_registers_1_5_Re : _GEN_1847; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1849 = 5'h6 == _GEN_1818 ? input_delay_registers_1_6_Re : _GEN_1848; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1850 = 5'h7 == _GEN_1818 ? input_delay_registers_1_7_Re : _GEN_1849; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1851 = 5'h8 == _GEN_1818 ? input_delay_registers_1_8_Re : _GEN_1850; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1852 = 5'h9 == _GEN_1818 ? input_delay_registers_1_9_Re : _GEN_1851; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1853 = 5'ha == _GEN_1818 ? input_delay_registers_1_10_Re : _GEN_1852; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1854 = 5'hb == _GEN_1818 ? input_delay_registers_1_11_Re : _GEN_1853; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1855 = 5'hc == _GEN_1818 ? input_delay_registers_1_12_Re : _GEN_1854; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1856 = 5'hd == _GEN_1818 ? input_delay_registers_1_13_Re : _GEN_1855; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1857 = 5'he == _GEN_1818 ? input_delay_registers_1_14_Re : _GEN_1856; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1858 = 5'hf == _GEN_1818 ? input_delay_registers_1_15_Re : _GEN_1857; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1859 = 5'h10 == _GEN_1818 ? input_delay_registers_1_16_Re : _GEN_1858; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1860 = 5'h11 == _GEN_1818 ? input_delay_registers_1_17_Re : _GEN_1859; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1861 = 5'h12 == _GEN_1818 ? input_delay_registers_1_18_Re : _GEN_1860; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1862 = 5'h13 == _GEN_1818 ? input_delay_registers_1_19_Re : _GEN_1861; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1863 = 5'h14 == _GEN_1818 ? input_delay_registers_1_20_Re : _GEN_1862; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1864 = 5'h15 == _GEN_1818 ? input_delay_registers_1_21_Re : _GEN_1863; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1865 = 5'h16 == _GEN_1818 ? input_delay_registers_1_22_Re : _GEN_1864; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1866 = 5'h17 == _GEN_1818 ? input_delay_registers_1_23_Re : _GEN_1865; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1876 = 2'h1 == cnt ? 5'h17 : 5'h0; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1877 = 2'h2 == cnt ? 5'h0 : _GEN_1876; // @[FFTDesigns.scala 2979:{32,32}]
  wire [4:0] _GEN_1878 = 2'h3 == cnt ? 5'h17 : _GEN_1877; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1880 = 5'h1 == _GEN_1878 ? input_delay_registers_1_1_Im : input_delay_registers_1_0_Im; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1881 = 5'h2 == _GEN_1878 ? input_delay_registers_1_2_Im : _GEN_1880; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1882 = 5'h3 == _GEN_1878 ? input_delay_registers_1_3_Im : _GEN_1881; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1883 = 5'h4 == _GEN_1878 ? input_delay_registers_1_4_Im : _GEN_1882; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1884 = 5'h5 == _GEN_1878 ? input_delay_registers_1_5_Im : _GEN_1883; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1885 = 5'h6 == _GEN_1878 ? input_delay_registers_1_6_Im : _GEN_1884; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1886 = 5'h7 == _GEN_1878 ? input_delay_registers_1_7_Im : _GEN_1885; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1887 = 5'h8 == _GEN_1878 ? input_delay_registers_1_8_Im : _GEN_1886; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1888 = 5'h9 == _GEN_1878 ? input_delay_registers_1_9_Im : _GEN_1887; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1889 = 5'ha == _GEN_1878 ? input_delay_registers_1_10_Im : _GEN_1888; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1890 = 5'hb == _GEN_1878 ? input_delay_registers_1_11_Im : _GEN_1889; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1891 = 5'hc == _GEN_1878 ? input_delay_registers_1_12_Im : _GEN_1890; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1892 = 5'hd == _GEN_1878 ? input_delay_registers_1_13_Im : _GEN_1891; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1893 = 5'he == _GEN_1878 ? input_delay_registers_1_14_Im : _GEN_1892; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1894 = 5'hf == _GEN_1878 ? input_delay_registers_1_15_Im : _GEN_1893; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1895 = 5'h10 == _GEN_1878 ? input_delay_registers_1_16_Im : _GEN_1894; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1896 = 5'h11 == _GEN_1878 ? input_delay_registers_1_17_Im : _GEN_1895; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1897 = 5'h12 == _GEN_1878 ? input_delay_registers_1_18_Im : _GEN_1896; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1898 = 5'h13 == _GEN_1878 ? input_delay_registers_1_19_Im : _GEN_1897; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1899 = 5'h14 == _GEN_1878 ? input_delay_registers_1_20_Im : _GEN_1898; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1900 = 5'h15 == _GEN_1878 ? input_delay_registers_1_21_Im : _GEN_1899; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1901 = 5'h16 == _GEN_1878 ? input_delay_registers_1_22_Im : _GEN_1900; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1902 = 5'h17 == _GEN_1878 ? input_delay_registers_1_23_Im : _GEN_1901; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1904 = 5'h1 == _GEN_1878 ? input_delay_registers_1_1_Re : input_delay_registers_1_0_Re; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1905 = 5'h2 == _GEN_1878 ? input_delay_registers_1_2_Re : _GEN_1904; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1906 = 5'h3 == _GEN_1878 ? input_delay_registers_1_3_Re : _GEN_1905; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1907 = 5'h4 == _GEN_1878 ? input_delay_registers_1_4_Re : _GEN_1906; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1908 = 5'h5 == _GEN_1878 ? input_delay_registers_1_5_Re : _GEN_1907; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1909 = 5'h6 == _GEN_1878 ? input_delay_registers_1_6_Re : _GEN_1908; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1910 = 5'h7 == _GEN_1878 ? input_delay_registers_1_7_Re : _GEN_1909; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1911 = 5'h8 == _GEN_1878 ? input_delay_registers_1_8_Re : _GEN_1910; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1912 = 5'h9 == _GEN_1878 ? input_delay_registers_1_9_Re : _GEN_1911; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1913 = 5'ha == _GEN_1878 ? input_delay_registers_1_10_Re : _GEN_1912; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1914 = 5'hb == _GEN_1878 ? input_delay_registers_1_11_Re : _GEN_1913; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1915 = 5'hc == _GEN_1878 ? input_delay_registers_1_12_Re : _GEN_1914; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1916 = 5'hd == _GEN_1878 ? input_delay_registers_1_13_Re : _GEN_1915; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1917 = 5'he == _GEN_1878 ? input_delay_registers_1_14_Re : _GEN_1916; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1918 = 5'hf == _GEN_1878 ? input_delay_registers_1_15_Re : _GEN_1917; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1919 = 5'h10 == _GEN_1878 ? input_delay_registers_1_16_Re : _GEN_1918; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1920 = 5'h11 == _GEN_1878 ? input_delay_registers_1_17_Re : _GEN_1919; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1921 = 5'h12 == _GEN_1878 ? input_delay_registers_1_18_Re : _GEN_1920; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1922 = 5'h13 == _GEN_1878 ? input_delay_registers_1_19_Re : _GEN_1921; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1923 = 5'h14 == _GEN_1878 ? input_delay_registers_1_20_Re : _GEN_1922; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1924 = 5'h15 == _GEN_1878 ? input_delay_registers_1_21_Re : _GEN_1923; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1925 = 5'h16 == _GEN_1878 ? input_delay_registers_1_22_Re : _GEN_1924; // @[FFTDesigns.scala 2979:{32,32}]
  wire [31:0] _GEN_1926 = 5'h17 == _GEN_1878 ? input_delay_registers_1_23_Re : _GEN_1925; // @[FFTDesigns.scala 2979:{32,32}]
  RAM_Block_mw RAM_Block_mw ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_clock),
    .io_in_raddr(RAM_Block_mw_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_io_in_data_1_Im),
    .io_re(RAM_Block_mw_io_re),
    .io_wr_0(RAM_Block_mw_io_wr_0),
    .io_wr_1(RAM_Block_mw_io_wr_1),
    .io_en(RAM_Block_mw_io_en),
    .io_out_data_Re(RAM_Block_mw_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_1 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_1_clock),
    .io_in_raddr(RAM_Block_mw_1_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_1_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_1_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_1_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_1_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_1_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_1_io_in_data_1_Im),
    .io_re(RAM_Block_mw_1_io_re),
    .io_wr_0(RAM_Block_mw_1_io_wr_0),
    .io_wr_1(RAM_Block_mw_1_io_wr_1),
    .io_en(RAM_Block_mw_1_io_en),
    .io_out_data_Re(RAM_Block_mw_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_1_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_2 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_2_clock),
    .io_in_raddr(RAM_Block_mw_2_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_2_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_2_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_2_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_2_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_2_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_2_io_in_data_1_Im),
    .io_re(RAM_Block_mw_2_io_re),
    .io_wr_0(RAM_Block_mw_2_io_wr_0),
    .io_wr_1(RAM_Block_mw_2_io_wr_1),
    .io_en(RAM_Block_mw_2_io_en),
    .io_out_data_Re(RAM_Block_mw_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_2_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_3 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_3_clock),
    .io_in_raddr(RAM_Block_mw_3_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_3_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_3_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_3_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_3_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_3_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_3_io_in_data_1_Im),
    .io_re(RAM_Block_mw_3_io_re),
    .io_wr_0(RAM_Block_mw_3_io_wr_0),
    .io_wr_1(RAM_Block_mw_3_io_wr_1),
    .io_en(RAM_Block_mw_3_io_en),
    .io_out_data_Re(RAM_Block_mw_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_3_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_4 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_4_clock),
    .io_in_raddr(RAM_Block_mw_4_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_4_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_4_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_4_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_4_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_4_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_4_io_in_data_1_Im),
    .io_re(RAM_Block_mw_4_io_re),
    .io_wr_0(RAM_Block_mw_4_io_wr_0),
    .io_wr_1(RAM_Block_mw_4_io_wr_1),
    .io_en(RAM_Block_mw_4_io_en),
    .io_out_data_Re(RAM_Block_mw_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_4_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_5 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_5_clock),
    .io_in_raddr(RAM_Block_mw_5_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_5_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_5_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_5_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_5_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_5_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_5_io_in_data_1_Im),
    .io_re(RAM_Block_mw_5_io_re),
    .io_wr_0(RAM_Block_mw_5_io_wr_0),
    .io_wr_1(RAM_Block_mw_5_io_wr_1),
    .io_en(RAM_Block_mw_5_io_en),
    .io_out_data_Re(RAM_Block_mw_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_5_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_6 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_6_clock),
    .io_in_raddr(RAM_Block_mw_6_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_6_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_6_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_6_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_6_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_6_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_6_io_in_data_1_Im),
    .io_re(RAM_Block_mw_6_io_re),
    .io_wr_0(RAM_Block_mw_6_io_wr_0),
    .io_wr_1(RAM_Block_mw_6_io_wr_1),
    .io_en(RAM_Block_mw_6_io_en),
    .io_out_data_Re(RAM_Block_mw_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_6_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_7 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_7_clock),
    .io_in_raddr(RAM_Block_mw_7_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_7_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_7_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_7_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_7_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_7_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_7_io_in_data_1_Im),
    .io_re(RAM_Block_mw_7_io_re),
    .io_wr_0(RAM_Block_mw_7_io_wr_0),
    .io_wr_1(RAM_Block_mw_7_io_wr_1),
    .io_en(RAM_Block_mw_7_io_en),
    .io_out_data_Re(RAM_Block_mw_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_7_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_8 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_8_clock),
    .io_in_raddr(RAM_Block_mw_8_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_8_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_8_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_8_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_8_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_8_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_8_io_in_data_1_Im),
    .io_re(RAM_Block_mw_8_io_re),
    .io_wr_0(RAM_Block_mw_8_io_wr_0),
    .io_wr_1(RAM_Block_mw_8_io_wr_1),
    .io_en(RAM_Block_mw_8_io_en),
    .io_out_data_Re(RAM_Block_mw_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_8_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_9 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_9_clock),
    .io_in_raddr(RAM_Block_mw_9_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_9_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_9_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_9_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_9_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_9_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_9_io_in_data_1_Im),
    .io_re(RAM_Block_mw_9_io_re),
    .io_wr_0(RAM_Block_mw_9_io_wr_0),
    .io_wr_1(RAM_Block_mw_9_io_wr_1),
    .io_en(RAM_Block_mw_9_io_en),
    .io_out_data_Re(RAM_Block_mw_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_9_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_10 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_10_clock),
    .io_in_raddr(RAM_Block_mw_10_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_10_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_10_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_10_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_10_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_10_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_10_io_in_data_1_Im),
    .io_re(RAM_Block_mw_10_io_re),
    .io_wr_0(RAM_Block_mw_10_io_wr_0),
    .io_wr_1(RAM_Block_mw_10_io_wr_1),
    .io_en(RAM_Block_mw_10_io_en),
    .io_out_data_Re(RAM_Block_mw_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_10_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_11 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_11_clock),
    .io_in_raddr(RAM_Block_mw_11_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_11_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_11_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_11_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_11_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_11_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_11_io_in_data_1_Im),
    .io_re(RAM_Block_mw_11_io_re),
    .io_wr_0(RAM_Block_mw_11_io_wr_0),
    .io_wr_1(RAM_Block_mw_11_io_wr_1),
    .io_en(RAM_Block_mw_11_io_en),
    .io_out_data_Re(RAM_Block_mw_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_11_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_12 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_12_clock),
    .io_in_raddr(RAM_Block_mw_12_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_12_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_12_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_12_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_12_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_12_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_12_io_in_data_1_Im),
    .io_re(RAM_Block_mw_12_io_re),
    .io_wr_0(RAM_Block_mw_12_io_wr_0),
    .io_wr_1(RAM_Block_mw_12_io_wr_1),
    .io_en(RAM_Block_mw_12_io_en),
    .io_out_data_Re(RAM_Block_mw_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_12_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_13 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_13_clock),
    .io_in_raddr(RAM_Block_mw_13_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_13_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_13_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_13_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_13_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_13_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_13_io_in_data_1_Im),
    .io_re(RAM_Block_mw_13_io_re),
    .io_wr_0(RAM_Block_mw_13_io_wr_0),
    .io_wr_1(RAM_Block_mw_13_io_wr_1),
    .io_en(RAM_Block_mw_13_io_en),
    .io_out_data_Re(RAM_Block_mw_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_13_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_14 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_14_clock),
    .io_in_raddr(RAM_Block_mw_14_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_14_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_14_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_14_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_14_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_14_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_14_io_in_data_1_Im),
    .io_re(RAM_Block_mw_14_io_re),
    .io_wr_0(RAM_Block_mw_14_io_wr_0),
    .io_wr_1(RAM_Block_mw_14_io_wr_1),
    .io_en(RAM_Block_mw_14_io_en),
    .io_out_data_Re(RAM_Block_mw_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_14_io_out_data_Im)
  );
  RAM_Block_mw RAM_Block_mw_15 ( // @[FFTDesigns.scala 2837:26]
    .clock(RAM_Block_mw_15_clock),
    .io_in_raddr(RAM_Block_mw_15_io_in_raddr),
    .io_in_waddr_0(RAM_Block_mw_15_io_in_waddr_0),
    .io_in_waddr_1(RAM_Block_mw_15_io_in_waddr_1),
    .io_in_data_0_Re(RAM_Block_mw_15_io_in_data_0_Re),
    .io_in_data_0_Im(RAM_Block_mw_15_io_in_data_0_Im),
    .io_in_data_1_Re(RAM_Block_mw_15_io_in_data_1_Re),
    .io_in_data_1_Im(RAM_Block_mw_15_io_in_data_1_Im),
    .io_re(RAM_Block_mw_15_io_re),
    .io_wr_0(RAM_Block_mw_15_io_wr_0),
    .io_wr_1(RAM_Block_mw_15_io_wr_1),
    .io_en(RAM_Block_mw_15_io_en),
    .io_out_data_Re(RAM_Block_mw_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_mw_15_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_clock),
    .io_in_raddr(RAM_Block_io_in_raddr),
    .io_in_waddr(RAM_Block_io_in_waddr),
    .io_in_data_Re(RAM_Block_io_in_data_Re),
    .io_in_data_Im(RAM_Block_io_in_data_Im),
    .io_re(RAM_Block_io_re),
    .io_wr(RAM_Block_io_wr),
    .io_en(RAM_Block_io_en),
    .io_out_data_Re(RAM_Block_io_out_data_Re),
    .io_out_data_Im(RAM_Block_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_1 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_1_clock),
    .io_in_raddr(RAM_Block_1_io_in_raddr),
    .io_in_waddr(RAM_Block_1_io_in_waddr),
    .io_in_data_Re(RAM_Block_1_io_in_data_Re),
    .io_in_data_Im(RAM_Block_1_io_in_data_Im),
    .io_re(RAM_Block_1_io_re),
    .io_wr(RAM_Block_1_io_wr),
    .io_en(RAM_Block_1_io_en),
    .io_out_data_Re(RAM_Block_1_io_out_data_Re),
    .io_out_data_Im(RAM_Block_1_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_2 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_2_clock),
    .io_in_raddr(RAM_Block_2_io_in_raddr),
    .io_in_waddr(RAM_Block_2_io_in_waddr),
    .io_in_data_Re(RAM_Block_2_io_in_data_Re),
    .io_in_data_Im(RAM_Block_2_io_in_data_Im),
    .io_re(RAM_Block_2_io_re),
    .io_wr(RAM_Block_2_io_wr),
    .io_en(RAM_Block_2_io_en),
    .io_out_data_Re(RAM_Block_2_io_out_data_Re),
    .io_out_data_Im(RAM_Block_2_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_3 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_3_clock),
    .io_in_raddr(RAM_Block_3_io_in_raddr),
    .io_in_waddr(RAM_Block_3_io_in_waddr),
    .io_in_data_Re(RAM_Block_3_io_in_data_Re),
    .io_in_data_Im(RAM_Block_3_io_in_data_Im),
    .io_re(RAM_Block_3_io_re),
    .io_wr(RAM_Block_3_io_wr),
    .io_en(RAM_Block_3_io_en),
    .io_out_data_Re(RAM_Block_3_io_out_data_Re),
    .io_out_data_Im(RAM_Block_3_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_4 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_4_clock),
    .io_in_raddr(RAM_Block_4_io_in_raddr),
    .io_in_waddr(RAM_Block_4_io_in_waddr),
    .io_in_data_Re(RAM_Block_4_io_in_data_Re),
    .io_in_data_Im(RAM_Block_4_io_in_data_Im),
    .io_re(RAM_Block_4_io_re),
    .io_wr(RAM_Block_4_io_wr),
    .io_en(RAM_Block_4_io_en),
    .io_out_data_Re(RAM_Block_4_io_out_data_Re),
    .io_out_data_Im(RAM_Block_4_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_5 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_5_clock),
    .io_in_raddr(RAM_Block_5_io_in_raddr),
    .io_in_waddr(RAM_Block_5_io_in_waddr),
    .io_in_data_Re(RAM_Block_5_io_in_data_Re),
    .io_in_data_Im(RAM_Block_5_io_in_data_Im),
    .io_re(RAM_Block_5_io_re),
    .io_wr(RAM_Block_5_io_wr),
    .io_en(RAM_Block_5_io_en),
    .io_out_data_Re(RAM_Block_5_io_out_data_Re),
    .io_out_data_Im(RAM_Block_5_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_6 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_6_clock),
    .io_in_raddr(RAM_Block_6_io_in_raddr),
    .io_in_waddr(RAM_Block_6_io_in_waddr),
    .io_in_data_Re(RAM_Block_6_io_in_data_Re),
    .io_in_data_Im(RAM_Block_6_io_in_data_Im),
    .io_re(RAM_Block_6_io_re),
    .io_wr(RAM_Block_6_io_wr),
    .io_en(RAM_Block_6_io_en),
    .io_out_data_Re(RAM_Block_6_io_out_data_Re),
    .io_out_data_Im(RAM_Block_6_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_7 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_7_clock),
    .io_in_raddr(RAM_Block_7_io_in_raddr),
    .io_in_waddr(RAM_Block_7_io_in_waddr),
    .io_in_data_Re(RAM_Block_7_io_in_data_Re),
    .io_in_data_Im(RAM_Block_7_io_in_data_Im),
    .io_re(RAM_Block_7_io_re),
    .io_wr(RAM_Block_7_io_wr),
    .io_en(RAM_Block_7_io_en),
    .io_out_data_Re(RAM_Block_7_io_out_data_Re),
    .io_out_data_Im(RAM_Block_7_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_8 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_8_clock),
    .io_in_raddr(RAM_Block_8_io_in_raddr),
    .io_in_waddr(RAM_Block_8_io_in_waddr),
    .io_in_data_Re(RAM_Block_8_io_in_data_Re),
    .io_in_data_Im(RAM_Block_8_io_in_data_Im),
    .io_re(RAM_Block_8_io_re),
    .io_wr(RAM_Block_8_io_wr),
    .io_en(RAM_Block_8_io_en),
    .io_out_data_Re(RAM_Block_8_io_out_data_Re),
    .io_out_data_Im(RAM_Block_8_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_9 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_9_clock),
    .io_in_raddr(RAM_Block_9_io_in_raddr),
    .io_in_waddr(RAM_Block_9_io_in_waddr),
    .io_in_data_Re(RAM_Block_9_io_in_data_Re),
    .io_in_data_Im(RAM_Block_9_io_in_data_Im),
    .io_re(RAM_Block_9_io_re),
    .io_wr(RAM_Block_9_io_wr),
    .io_en(RAM_Block_9_io_en),
    .io_out_data_Re(RAM_Block_9_io_out_data_Re),
    .io_out_data_Im(RAM_Block_9_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_10 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_10_clock),
    .io_in_raddr(RAM_Block_10_io_in_raddr),
    .io_in_waddr(RAM_Block_10_io_in_waddr),
    .io_in_data_Re(RAM_Block_10_io_in_data_Re),
    .io_in_data_Im(RAM_Block_10_io_in_data_Im),
    .io_re(RAM_Block_10_io_re),
    .io_wr(RAM_Block_10_io_wr),
    .io_en(RAM_Block_10_io_en),
    .io_out_data_Re(RAM_Block_10_io_out_data_Re),
    .io_out_data_Im(RAM_Block_10_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_11 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_11_clock),
    .io_in_raddr(RAM_Block_11_io_in_raddr),
    .io_in_waddr(RAM_Block_11_io_in_waddr),
    .io_in_data_Re(RAM_Block_11_io_in_data_Re),
    .io_in_data_Im(RAM_Block_11_io_in_data_Im),
    .io_re(RAM_Block_11_io_re),
    .io_wr(RAM_Block_11_io_wr),
    .io_en(RAM_Block_11_io_en),
    .io_out_data_Re(RAM_Block_11_io_out_data_Re),
    .io_out_data_Im(RAM_Block_11_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_12 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_12_clock),
    .io_in_raddr(RAM_Block_12_io_in_raddr),
    .io_in_waddr(RAM_Block_12_io_in_waddr),
    .io_in_data_Re(RAM_Block_12_io_in_data_Re),
    .io_in_data_Im(RAM_Block_12_io_in_data_Im),
    .io_re(RAM_Block_12_io_re),
    .io_wr(RAM_Block_12_io_wr),
    .io_en(RAM_Block_12_io_en),
    .io_out_data_Re(RAM_Block_12_io_out_data_Re),
    .io_out_data_Im(RAM_Block_12_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_13 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_13_clock),
    .io_in_raddr(RAM_Block_13_io_in_raddr),
    .io_in_waddr(RAM_Block_13_io_in_waddr),
    .io_in_data_Re(RAM_Block_13_io_in_data_Re),
    .io_in_data_Im(RAM_Block_13_io_in_data_Im),
    .io_re(RAM_Block_13_io_re),
    .io_wr(RAM_Block_13_io_wr),
    .io_en(RAM_Block_13_io_en),
    .io_out_data_Re(RAM_Block_13_io_out_data_Re),
    .io_out_data_Im(RAM_Block_13_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_14 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_14_clock),
    .io_in_raddr(RAM_Block_14_io_in_raddr),
    .io_in_waddr(RAM_Block_14_io_in_waddr),
    .io_in_data_Re(RAM_Block_14_io_in_data_Re),
    .io_in_data_Im(RAM_Block_14_io_in_data_Im),
    .io_re(RAM_Block_14_io_re),
    .io_wr(RAM_Block_14_io_wr),
    .io_en(RAM_Block_14_io_en),
    .io_out_data_Re(RAM_Block_14_io_out_data_Re),
    .io_out_data_Im(RAM_Block_14_io_out_data_Im)
  );
  RAM_Block_192 RAM_Block_15 ( // @[FFTDesigns.scala 2841:26]
    .clock(RAM_Block_15_clock),
    .io_in_raddr(RAM_Block_15_io_in_raddr),
    .io_in_waddr(RAM_Block_15_io_in_waddr),
    .io_in_data_Re(RAM_Block_15_io_in_data_Re),
    .io_in_data_Im(RAM_Block_15_io_in_data_Im),
    .io_re(RAM_Block_15_io_re),
    .io_wr(RAM_Block_15_io_wr),
    .io_en(RAM_Block_15_io_en),
    .io_out_data_Re(RAM_Block_15_io_out_data_Re),
    .io_out_data_Im(RAM_Block_15_io_out_data_Im)
  );
  PermutationModuleStreamed PermutationModuleStreamed ( // @[FFTDesigns.scala 2907:28]
    .io_in_0_Re(PermutationModuleStreamed_io_in_0_Re),
    .io_in_0_Im(PermutationModuleStreamed_io_in_0_Im),
    .io_in_1_Re(PermutationModuleStreamed_io_in_1_Re),
    .io_in_1_Im(PermutationModuleStreamed_io_in_1_Im),
    .io_in_2_Re(PermutationModuleStreamed_io_in_2_Re),
    .io_in_2_Im(PermutationModuleStreamed_io_in_2_Im),
    .io_in_3_Re(PermutationModuleStreamed_io_in_3_Re),
    .io_in_3_Im(PermutationModuleStreamed_io_in_3_Im),
    .io_in_4_Re(PermutationModuleStreamed_io_in_4_Re),
    .io_in_4_Im(PermutationModuleStreamed_io_in_4_Im),
    .io_in_5_Re(PermutationModuleStreamed_io_in_5_Re),
    .io_in_5_Im(PermutationModuleStreamed_io_in_5_Im),
    .io_in_6_Re(PermutationModuleStreamed_io_in_6_Re),
    .io_in_6_Im(PermutationModuleStreamed_io_in_6_Im),
    .io_in_7_Re(PermutationModuleStreamed_io_in_7_Re),
    .io_in_7_Im(PermutationModuleStreamed_io_in_7_Im),
    .io_in_8_Re(PermutationModuleStreamed_io_in_8_Re),
    .io_in_8_Im(PermutationModuleStreamed_io_in_8_Im),
    .io_in_9_Re(PermutationModuleStreamed_io_in_9_Re),
    .io_in_9_Im(PermutationModuleStreamed_io_in_9_Im),
    .io_in_10_Re(PermutationModuleStreamed_io_in_10_Re),
    .io_in_10_Im(PermutationModuleStreamed_io_in_10_Im),
    .io_in_11_Re(PermutationModuleStreamed_io_in_11_Re),
    .io_in_11_Im(PermutationModuleStreamed_io_in_11_Im),
    .io_in_12_Re(PermutationModuleStreamed_io_in_12_Re),
    .io_in_12_Im(PermutationModuleStreamed_io_in_12_Im),
    .io_in_13_Re(PermutationModuleStreamed_io_in_13_Re),
    .io_in_13_Im(PermutationModuleStreamed_io_in_13_Im),
    .io_in_14_Re(PermutationModuleStreamed_io_in_14_Re),
    .io_in_14_Im(PermutationModuleStreamed_io_in_14_Im),
    .io_in_15_Re(PermutationModuleStreamed_io_in_15_Re),
    .io_in_15_Im(PermutationModuleStreamed_io_in_15_Im),
    .io_in_config_0(PermutationModuleStreamed_io_in_config_0),
    .io_in_config_1(PermutationModuleStreamed_io_in_config_1),
    .io_in_config_2(PermutationModuleStreamed_io_in_config_2),
    .io_in_config_3(PermutationModuleStreamed_io_in_config_3),
    .io_in_config_4(PermutationModuleStreamed_io_in_config_4),
    .io_in_config_5(PermutationModuleStreamed_io_in_config_5),
    .io_in_config_6(PermutationModuleStreamed_io_in_config_6),
    .io_in_config_7(PermutationModuleStreamed_io_in_config_7),
    .io_in_config_8(PermutationModuleStreamed_io_in_config_8),
    .io_in_config_9(PermutationModuleStreamed_io_in_config_9),
    .io_in_config_10(PermutationModuleStreamed_io_in_config_10),
    .io_in_config_11(PermutationModuleStreamed_io_in_config_11),
    .io_in_config_12(PermutationModuleStreamed_io_in_config_12),
    .io_in_config_13(PermutationModuleStreamed_io_in_config_13),
    .io_in_config_14(PermutationModuleStreamed_io_in_config_14),
    .io_out_0_Re(PermutationModuleStreamed_io_out_0_Re),
    .io_out_0_Im(PermutationModuleStreamed_io_out_0_Im),
    .io_out_1_Re(PermutationModuleStreamed_io_out_1_Re),
    .io_out_1_Im(PermutationModuleStreamed_io_out_1_Im),
    .io_out_2_Re(PermutationModuleStreamed_io_out_2_Re),
    .io_out_2_Im(PermutationModuleStreamed_io_out_2_Im),
    .io_out_3_Re(PermutationModuleStreamed_io_out_3_Re),
    .io_out_3_Im(PermutationModuleStreamed_io_out_3_Im),
    .io_out_4_Re(PermutationModuleStreamed_io_out_4_Re),
    .io_out_4_Im(PermutationModuleStreamed_io_out_4_Im),
    .io_out_5_Re(PermutationModuleStreamed_io_out_5_Re),
    .io_out_5_Im(PermutationModuleStreamed_io_out_5_Im),
    .io_out_6_Re(PermutationModuleStreamed_io_out_6_Re),
    .io_out_6_Im(PermutationModuleStreamed_io_out_6_Im),
    .io_out_7_Re(PermutationModuleStreamed_io_out_7_Re),
    .io_out_7_Im(PermutationModuleStreamed_io_out_7_Im),
    .io_out_8_Re(PermutationModuleStreamed_io_out_8_Re),
    .io_out_8_Im(PermutationModuleStreamed_io_out_8_Im),
    .io_out_9_Re(PermutationModuleStreamed_io_out_9_Re),
    .io_out_9_Im(PermutationModuleStreamed_io_out_9_Im),
    .io_out_10_Re(PermutationModuleStreamed_io_out_10_Re),
    .io_out_10_Im(PermutationModuleStreamed_io_out_10_Im),
    .io_out_11_Re(PermutationModuleStreamed_io_out_11_Re),
    .io_out_11_Im(PermutationModuleStreamed_io_out_11_Im),
    .io_out_12_Re(PermutationModuleStreamed_io_out_12_Re),
    .io_out_12_Im(PermutationModuleStreamed_io_out_12_Im),
    .io_out_13_Re(PermutationModuleStreamed_io_out_13_Re),
    .io_out_13_Im(PermutationModuleStreamed_io_out_13_Im),
    .io_out_14_Re(PermutationModuleStreamed_io_out_14_Re),
    .io_out_14_Im(PermutationModuleStreamed_io_out_14_Im),
    .io_out_15_Re(PermutationModuleStreamed_io_out_15_Re),
    .io_out_15_Im(PermutationModuleStreamed_io_out_15_Im)
  );
  M0_Config_ROM_6 M0_Config_ROM ( // @[FFTDesigns.scala 2908:29]
    .io_in_cnt(M0_Config_ROM_io_in_cnt),
    .io_out_0(M0_Config_ROM_io_out_0),
    .io_out_1(M0_Config_ROM_io_out_1),
    .io_out_2(M0_Config_ROM_io_out_2),
    .io_out_3(M0_Config_ROM_io_out_3),
    .io_out_4(M0_Config_ROM_io_out_4),
    .io_out_5(M0_Config_ROM_io_out_5),
    .io_out_6(M0_Config_ROM_io_out_6),
    .io_out_7(M0_Config_ROM_io_out_7),
    .io_out_8(M0_Config_ROM_io_out_8),
    .io_out_9(M0_Config_ROM_io_out_9),
    .io_out_10(M0_Config_ROM_io_out_10),
    .io_out_11(M0_Config_ROM_io_out_11),
    .io_out_12(M0_Config_ROM_io_out_12),
    .io_out_13(M0_Config_ROM_io_out_13),
    .io_out_14(M0_Config_ROM_io_out_14),
    .io_out_15(M0_Config_ROM_io_out_15)
  );
  M1_Config_ROM_6 M1_Config_ROM ( // @[FFTDesigns.scala 2909:29]
    .io_in_cnt(M1_Config_ROM_io_in_cnt),
    .io_out_0(M1_Config_ROM_io_out_0),
    .io_out_1(M1_Config_ROM_io_out_1),
    .io_out_2(M1_Config_ROM_io_out_2),
    .io_out_3(M1_Config_ROM_io_out_3),
    .io_out_4(M1_Config_ROM_io_out_4),
    .io_out_5(M1_Config_ROM_io_out_5),
    .io_out_6(M1_Config_ROM_io_out_6),
    .io_out_7(M1_Config_ROM_io_out_7),
    .io_out_8(M1_Config_ROM_io_out_8),
    .io_out_9(M1_Config_ROM_io_out_9),
    .io_out_10(M1_Config_ROM_io_out_10),
    .io_out_11(M1_Config_ROM_io_out_11),
    .io_out_12(M1_Config_ROM_io_out_12),
    .io_out_13(M1_Config_ROM_io_out_13),
    .io_out_14(M1_Config_ROM_io_out_14),
    .io_out_15(M1_Config_ROM_io_out_15)
  );
  Streaming_Permute_Config_6 Streaming_Permute_Config ( // @[FFTDesigns.scala 2910:31]
    .io_in_cnt(Streaming_Permute_Config_io_in_cnt),
    .io_out_0(Streaming_Permute_Config_io_out_0),
    .io_out_1(Streaming_Permute_Config_io_out_1),
    .io_out_2(Streaming_Permute_Config_io_out_2),
    .io_out_3(Streaming_Permute_Config_io_out_3),
    .io_out_4(Streaming_Permute_Config_io_out_4),
    .io_out_5(Streaming_Permute_Config_io_out_5),
    .io_out_6(Streaming_Permute_Config_io_out_6),
    .io_out_7(Streaming_Permute_Config_io_out_7),
    .io_out_8(Streaming_Permute_Config_io_out_8),
    .io_out_9(Streaming_Permute_Config_io_out_9),
    .io_out_10(Streaming_Permute_Config_io_out_10),
    .io_out_11(Streaming_Permute_Config_io_out_11),
    .io_out_12(Streaming_Permute_Config_io_out_12),
    .io_out_13(Streaming_Permute_Config_io_out_13),
    .io_out_14(Streaming_Permute_Config_io_out_14)
  );
  assign io_out_0_Re = RAM_Block_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_0_Im = RAM_Block_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_1_Re = RAM_Block_1_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_1_Im = RAM_Block_1_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_2_Re = RAM_Block_2_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_2_Im = RAM_Block_2_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_3_Re = RAM_Block_3_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_3_Im = RAM_Block_3_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_4_Re = RAM_Block_4_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_4_Im = RAM_Block_4_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_5_Re = RAM_Block_5_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_5_Im = RAM_Block_5_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_6_Re = RAM_Block_6_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_6_Im = RAM_Block_6_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_7_Re = RAM_Block_7_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_7_Im = RAM_Block_7_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_8_Re = RAM_Block_8_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_8_Im = RAM_Block_8_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_9_Re = RAM_Block_9_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_9_Im = RAM_Block_9_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_10_Re = RAM_Block_10_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_10_Im = RAM_Block_10_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_11_Re = RAM_Block_11_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_11_Im = RAM_Block_11_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_12_Re = RAM_Block_12_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_12_Im = RAM_Block_12_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_13_Re = RAM_Block_13_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_13_Im = RAM_Block_13_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_14_Re = RAM_Block_14_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_14_Im = RAM_Block_14_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_15_Re = RAM_Block_15_io_out_data_Re; // @[FFTDesigns.scala 2840:{23,23}]
  assign io_out_15_Im = RAM_Block_15_io_out_data_Im; // @[FFTDesigns.scala 2840:{23,23}]
  assign RAM_Block_mw_clock = clock;
  assign RAM_Block_mw_io_in_raddr = M0_0_re ? _M0_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_io_in_data_0_Re = M0_0_re ? _GEN_66 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_io_in_data_0_Im = M0_0_re ? _GEN_42 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_io_in_data_1_Re = M0_0_re ? _GEN_126 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_io_in_data_1_Im = M0_0_re ? _GEN_102 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_io_wr_1 = M0_0_re & _GEN_70; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_1_clock = clock;
  assign RAM_Block_mw_1_io_in_raddr = M0_0_re ? _M0_1_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_1_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_1_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_1_io_in_data_0_Re = M0_0_re ? _GEN_186 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_1_io_in_data_0_Im = M0_0_re ? _GEN_162 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_1_io_in_data_1_Re = M0_0_re ? _GEN_246 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_1_io_in_data_1_Im = M0_0_re ? _GEN_222 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_1_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_1_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_1_io_wr_1 = M0_0_re & _GEN_70; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_1_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_2_clock = clock;
  assign RAM_Block_mw_2_io_in_raddr = M0_0_re ? _M0_2_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_2_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_2_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_2_io_in_data_0_Re = M0_0_re ? _GEN_306 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_2_io_in_data_0_Im = M0_0_re ? _GEN_282 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_2_io_in_data_1_Re = M0_0_re ? _GEN_366 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_2_io_in_data_1_Im = M0_0_re ? _GEN_342 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_2_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_2_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_2_io_wr_1 = M0_0_re & _GEN_70; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_2_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_3_clock = clock;
  assign RAM_Block_mw_3_io_in_raddr = M0_0_re ? _M0_3_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_3_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_3_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_3_io_in_data_0_Re = M0_0_re ? _GEN_426 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_3_io_in_data_0_Im = M0_0_re ? _GEN_402 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_3_io_in_data_1_Re = M0_0_re ? _GEN_486 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_3_io_in_data_1_Im = M0_0_re ? _GEN_462 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_3_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_3_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_3_io_wr_1 = M0_0_re & _GEN_70; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_3_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_4_clock = clock;
  assign RAM_Block_mw_4_io_in_raddr = M0_0_re ? _M0_4_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_4_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_4_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_4_io_in_data_0_Re = M0_0_re ? _GEN_546 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_4_io_in_data_0_Im = M0_0_re ? _GEN_522 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_4_io_in_data_1_Re = M0_0_re ? _GEN_606 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_4_io_in_data_1_Im = M0_0_re ? _GEN_582 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_4_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_4_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_4_io_wr_1 = M0_0_re & _GEN_70; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_4_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_5_clock = clock;
  assign RAM_Block_mw_5_io_in_raddr = M0_0_re ? _M0_5_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_5_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_5_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_5_io_in_data_0_Re = M0_0_re ? _GEN_666 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_5_io_in_data_0_Im = M0_0_re ? _GEN_642 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_5_io_in_data_1_Re = M0_0_re ? _GEN_726 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_5_io_in_data_1_Im = M0_0_re ? _GEN_702 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_5_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_5_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_5_io_wr_1 = M0_0_re & _GEN_70; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_5_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_6_clock = clock;
  assign RAM_Block_mw_6_io_in_raddr = M0_0_re ? _M0_6_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_6_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_6_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_6_io_in_data_0_Re = M0_0_re ? _GEN_786 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_6_io_in_data_0_Im = M0_0_re ? _GEN_762 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_6_io_in_data_1_Re = M0_0_re ? _GEN_846 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_6_io_in_data_1_Im = M0_0_re ? _GEN_822 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_6_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_6_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_6_io_wr_1 = M0_0_re & _GEN_70; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_6_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_7_clock = clock;
  assign RAM_Block_mw_7_io_in_raddr = M0_0_re ? _M0_7_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_7_io_in_waddr_0 = M0_0_re ? _M0_0_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_7_io_in_waddr_1 = M0_0_re ? _M0_0_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_7_io_in_data_0_Re = M0_0_re ? _GEN_906 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_7_io_in_data_0_Im = M0_0_re ? _GEN_882 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_7_io_in_data_1_Re = M0_0_re ? _GEN_966 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_7_io_in_data_1_Im = M0_0_re ? _GEN_942 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_7_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_7_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_7_io_wr_1 = M0_0_re & _GEN_70; // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_7_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_8_clock = clock;
  assign RAM_Block_mw_8_io_in_raddr = M0_0_re ? _M0_8_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_8_io_in_waddr_0 = M0_0_re ? _M0_8_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_8_io_in_waddr_1 = M0_0_re ? _M0_8_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_8_io_in_data_0_Re = M0_0_re ? _GEN_1026 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_8_io_in_data_0_Im = M0_0_re ? _GEN_1002 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_8_io_in_data_1_Re = M0_0_re ? _GEN_1086 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_8_io_in_data_1_Im = M0_0_re ? _GEN_1062 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_8_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_8_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_8_io_wr_1 = M0_0_re & (2'h3 == cnt | _GEN_1029); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_8_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_9_clock = clock;
  assign RAM_Block_mw_9_io_in_raddr = M0_0_re ? _M0_9_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_9_io_in_waddr_0 = M0_0_re ? _M0_8_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_9_io_in_waddr_1 = M0_0_re ? _M0_8_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_9_io_in_data_0_Re = M0_0_re ? _GEN_1146 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_9_io_in_data_0_Im = M0_0_re ? _GEN_1122 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_9_io_in_data_1_Re = M0_0_re ? _GEN_1206 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_9_io_in_data_1_Im = M0_0_re ? _GEN_1182 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_9_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_9_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_9_io_wr_1 = M0_0_re & (2'h3 == cnt | _GEN_1029); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_9_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_10_clock = clock;
  assign RAM_Block_mw_10_io_in_raddr = M0_0_re ? _M0_10_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_10_io_in_waddr_0 = M0_0_re ? _M0_8_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_10_io_in_waddr_1 = M0_0_re ? _M0_8_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_10_io_in_data_0_Re = M0_0_re ? _GEN_1266 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_10_io_in_data_0_Im = M0_0_re ? _GEN_1242 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_10_io_in_data_1_Re = M0_0_re ? _GEN_1326 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_10_io_in_data_1_Im = M0_0_re ? _GEN_1302 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_10_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_10_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_10_io_wr_1 = M0_0_re & (2'h3 == cnt | _GEN_1029); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_10_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_11_clock = clock;
  assign RAM_Block_mw_11_io_in_raddr = M0_0_re ? _M0_11_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_11_io_in_waddr_0 = M0_0_re ? _M0_8_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_11_io_in_waddr_1 = M0_0_re ? _M0_8_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_11_io_in_data_0_Re = M0_0_re ? _GEN_1386 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_11_io_in_data_0_Im = M0_0_re ? _GEN_1362 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_11_io_in_data_1_Re = M0_0_re ? _GEN_1446 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_11_io_in_data_1_Im = M0_0_re ? _GEN_1422 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_11_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_11_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_11_io_wr_1 = M0_0_re & (2'h3 == cnt | _GEN_1029); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_11_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_12_clock = clock;
  assign RAM_Block_mw_12_io_in_raddr = M0_0_re ? _M0_12_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_12_io_in_waddr_0 = M0_0_re ? _M0_8_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_12_io_in_waddr_1 = M0_0_re ? _M0_8_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_12_io_in_data_0_Re = M0_0_re ? _GEN_1506 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_12_io_in_data_0_Im = M0_0_re ? _GEN_1482 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_12_io_in_data_1_Re = M0_0_re ? _GEN_1566 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_12_io_in_data_1_Im = M0_0_re ? _GEN_1542 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_12_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_12_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_12_io_wr_1 = M0_0_re & (2'h3 == cnt | _GEN_1029); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_12_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_13_clock = clock;
  assign RAM_Block_mw_13_io_in_raddr = M0_0_re ? _M0_13_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_13_io_in_waddr_0 = M0_0_re ? _M0_8_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_13_io_in_waddr_1 = M0_0_re ? _M0_8_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_13_io_in_data_0_Re = M0_0_re ? _GEN_1626 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_13_io_in_data_0_Im = M0_0_re ? _GEN_1602 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_13_io_in_data_1_Re = M0_0_re ? _GEN_1686 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_13_io_in_data_1_Im = M0_0_re ? _GEN_1662 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_13_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_13_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_13_io_wr_1 = M0_0_re & (2'h3 == cnt | _GEN_1029); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_13_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_14_clock = clock;
  assign RAM_Block_mw_14_io_in_raddr = M0_0_re ? _M0_14_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_14_io_in_waddr_0 = M0_0_re ? _M0_8_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_14_io_in_waddr_1 = M0_0_re ? _M0_8_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_14_io_in_data_0_Re = M0_0_re ? _GEN_1746 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_14_io_in_data_0_Im = M0_0_re ? _GEN_1722 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_14_io_in_data_1_Re = M0_0_re ? _GEN_1806 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_14_io_in_data_1_Im = M0_0_re ? _GEN_1782 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_14_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_14_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_14_io_wr_1 = M0_0_re & (2'h3 == cnt | _GEN_1029); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_14_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_15_clock = clock;
  assign RAM_Block_mw_15_io_in_raddr = M0_0_re ? _M0_15_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2950:26 3005:26]
  assign RAM_Block_mw_15_io_in_waddr_0 = M0_0_re ? _M0_8_in_waddr_0_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_15_io_in_waddr_1 = M0_0_re ? _M0_8_in_waddr_1_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2978:33 3006:26]
  assign RAM_Block_mw_15_io_in_data_0_Re = M0_0_re ? _GEN_1866 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_15_io_in_data_0_Im = M0_0_re ? _GEN_1842 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_15_io_in_data_1_Re = M0_0_re ? _GEN_1926 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_15_io_in_data_1_Im = M0_0_re ? _GEN_1902 : 32'h0; // @[FFTDesigns.scala 2914:33 2979:32 3007:25]
  assign RAM_Block_mw_15_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_15_io_wr_0 = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_mw_15_io_wr_1 = M0_0_re & (2'h3 == cnt | _GEN_1029); // @[FFTDesigns.scala 2914:33 2977:27 3001:20]
  assign RAM_Block_mw_15_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_clock = clock;
  assign RAM_Block_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_io_in_waddr = M0_0_re ? _M1_0_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_io_in_data_Re = PermutationModuleStreamed_io_out_0_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_io_in_data_Im = PermutationModuleStreamed_io_out_0_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_1_clock = clock;
  assign RAM_Block_1_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_1_io_in_waddr = M0_0_re ? _M1_1_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_1_io_in_data_Re = PermutationModuleStreamed_io_out_1_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_1_io_in_data_Im = PermutationModuleStreamed_io_out_1_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_1_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_1_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_1_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_2_clock = clock;
  assign RAM_Block_2_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_2_io_in_waddr = M0_0_re ? _M1_2_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_2_io_in_data_Re = PermutationModuleStreamed_io_out_2_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_2_io_in_data_Im = PermutationModuleStreamed_io_out_2_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_2_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_2_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_2_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_3_clock = clock;
  assign RAM_Block_3_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_3_io_in_waddr = M0_0_re ? _M1_3_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_3_io_in_data_Re = PermutationModuleStreamed_io_out_3_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_3_io_in_data_Im = PermutationModuleStreamed_io_out_3_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_3_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_3_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_3_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_4_clock = clock;
  assign RAM_Block_4_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_4_io_in_waddr = M0_0_re ? _M1_4_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_4_io_in_data_Re = PermutationModuleStreamed_io_out_4_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_4_io_in_data_Im = PermutationModuleStreamed_io_out_4_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_4_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_4_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_4_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_5_clock = clock;
  assign RAM_Block_5_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_5_io_in_waddr = M0_0_re ? _M1_5_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_5_io_in_data_Re = PermutationModuleStreamed_io_out_5_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_5_io_in_data_Im = PermutationModuleStreamed_io_out_5_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_5_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_5_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_5_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_6_clock = clock;
  assign RAM_Block_6_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_6_io_in_waddr = M0_0_re ? _M1_6_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_6_io_in_data_Re = PermutationModuleStreamed_io_out_6_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_6_io_in_data_Im = PermutationModuleStreamed_io_out_6_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_6_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_6_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_6_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_7_clock = clock;
  assign RAM_Block_7_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_7_io_in_waddr = M0_0_re ? _M1_7_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_7_io_in_data_Re = PermutationModuleStreamed_io_out_7_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_7_io_in_data_Im = PermutationModuleStreamed_io_out_7_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_7_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_7_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_7_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_8_clock = clock;
  assign RAM_Block_8_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_8_io_in_waddr = M0_0_re ? _M1_8_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_8_io_in_data_Re = PermutationModuleStreamed_io_out_8_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_8_io_in_data_Im = PermutationModuleStreamed_io_out_8_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_8_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_8_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_8_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_9_clock = clock;
  assign RAM_Block_9_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_9_io_in_waddr = M0_0_re ? _M1_9_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_9_io_in_data_Re = PermutationModuleStreamed_io_out_9_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_9_io_in_data_Im = PermutationModuleStreamed_io_out_9_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_9_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_9_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_9_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_10_clock = clock;
  assign RAM_Block_10_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_10_io_in_waddr = M0_0_re ? _M1_10_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_10_io_in_data_Re = PermutationModuleStreamed_io_out_10_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_10_io_in_data_Im = PermutationModuleStreamed_io_out_10_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_10_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_10_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_10_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_11_clock = clock;
  assign RAM_Block_11_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_11_io_in_waddr = M0_0_re ? _M1_11_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_11_io_in_data_Re = PermutationModuleStreamed_io_out_11_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_11_io_in_data_Im = PermutationModuleStreamed_io_out_11_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_11_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_11_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_11_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_12_clock = clock;
  assign RAM_Block_12_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_12_io_in_waddr = M0_0_re ? _M1_12_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_12_io_in_data_Re = PermutationModuleStreamed_io_out_12_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_12_io_in_data_Im = PermutationModuleStreamed_io_out_12_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_12_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_12_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_12_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_13_clock = clock;
  assign RAM_Block_13_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_13_io_in_waddr = M0_0_re ? _M1_13_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_13_io_in_data_Re = PermutationModuleStreamed_io_out_13_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_13_io_in_data_Im = PermutationModuleStreamed_io_out_13_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_13_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_13_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_13_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_14_clock = clock;
  assign RAM_Block_14_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_14_io_in_waddr = M0_0_re ? _M1_14_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_14_io_in_data_Re = PermutationModuleStreamed_io_out_14_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_14_io_in_data_Im = PermutationModuleStreamed_io_out_14_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_14_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_14_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_14_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_15_clock = clock;
  assign RAM_Block_15_io_in_raddr = M0_0_re ? _M1_0_in_raddr_T_3 : 4'h0; // @[FFTDesigns.scala 2914:33 2951:26 3008:26]
  assign RAM_Block_15_io_in_waddr = M0_0_re ? _M1_15_in_waddr_T_2 : 4'h0; // @[FFTDesigns.scala 2914:33 2952:26 3009:26]
  assign RAM_Block_15_io_in_data_Re = PermutationModuleStreamed_io_out_15_Re; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_15_io_in_data_Im = PermutationModuleStreamed_io_out_15_Im; // @[FFTDesigns.scala 2914:33 2953:25 3010:25]
  assign RAM_Block_15_io_re = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_15_io_wr = |_T; // @[FFTDesigns.scala 2914:28]
  assign RAM_Block_15_io_en = |_T; // @[FFTDesigns.scala 2914:28]
  assign PermutationModuleStreamed_io_in_0_Re = RAM_Block_mw_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_0_Im = RAM_Block_mw_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_1_Re = RAM_Block_mw_1_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_1_Im = RAM_Block_mw_1_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_2_Re = RAM_Block_mw_2_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_2_Im = RAM_Block_mw_2_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_3_Re = RAM_Block_mw_3_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_3_Im = RAM_Block_mw_3_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_4_Re = RAM_Block_mw_4_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_4_Im = RAM_Block_mw_4_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_5_Re = RAM_Block_mw_5_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_5_Im = RAM_Block_mw_5_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_6_Re = RAM_Block_mw_6_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_6_Im = RAM_Block_mw_6_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_7_Re = RAM_Block_mw_7_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_7_Im = RAM_Block_mw_7_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_8_Re = RAM_Block_mw_8_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_8_Im = RAM_Block_mw_8_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_9_Re = RAM_Block_mw_9_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_9_Im = RAM_Block_mw_9_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_10_Re = RAM_Block_mw_10_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_10_Im = RAM_Block_mw_10_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_11_Re = RAM_Block_mw_11_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_11_Im = RAM_Block_mw_11_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_12_Re = RAM_Block_mw_12_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_12_Im = RAM_Block_mw_12_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_13_Re = RAM_Block_mw_13_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_13_Im = RAM_Block_mw_13_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_14_Re = RAM_Block_mw_14_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_14_Im = RAM_Block_mw_14_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_15_Re = RAM_Block_mw_15_io_out_data_Re; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_15_Im = RAM_Block_mw_15_io_out_data_Im; // @[FFTDesigns.scala 2836:{23,23}]
  assign PermutationModuleStreamed_io_in_config_0 = Streaming_Permute_Config_io_out_0; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_1 = Streaming_Permute_Config_io_out_1; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_2 = Streaming_Permute_Config_io_out_2; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_3 = Streaming_Permute_Config_io_out_3; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_4 = Streaming_Permute_Config_io_out_4; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_5 = Streaming_Permute_Config_io_out_5; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_6 = Streaming_Permute_Config_io_out_6; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_7 = Streaming_Permute_Config_io_out_7; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_8 = Streaming_Permute_Config_io_out_8; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_9 = Streaming_Permute_Config_io_out_9; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_10 = Streaming_Permute_Config_io_out_10; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_11 = Streaming_Permute_Config_io_out_11; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_12 = Streaming_Permute_Config_io_out_12; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_13 = Streaming_Permute_Config_io_out_13; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign PermutationModuleStreamed_io_in_config_14 = Streaming_Permute_Config_io_out_14; // @[FFTDesigns.scala 2914:33 2954:33 3011:33]
  assign M0_Config_ROM_io_in_cnt = cnt2; // @[FFTDesigns.scala 3021:24]
  assign M1_Config_ROM_io_in_cnt = cnt2; // @[FFTDesigns.scala 3022:24]
  assign Streaming_Permute_Config_io_in_cnt = cnt2; // @[FFTDesigns.scala 3023:26]
  always @(posedge clock) begin
    offset_switch <= M0_0_re & _GEN_6; // @[FFTDesigns.scala 2914:33 3017:23]
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_0_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_0_Re <= io_in_0_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_0_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_0_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_0_Im <= io_in_0_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_0_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_1_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_1_Re <= io_in_1_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_1_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_1_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_1_Im <= io_in_1_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_1_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_2_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_2_Re <= io_in_2_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_2_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_2_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_2_Im <= io_in_2_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_2_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_3_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_3_Re <= io_in_3_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_3_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_3_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_3_Im <= io_in_3_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_3_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_4_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_4_Re <= io_in_4_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_4_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_4_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_4_Im <= io_in_4_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_4_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_5_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_5_Re <= io_in_5_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_5_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_5_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_5_Im <= io_in_5_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_5_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_6_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_6_Re <= io_in_6_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_6_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_6_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_6_Im <= io_in_6_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_6_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_7_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_7_Re <= io_in_7_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_7_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_7_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_7_Im <= io_in_7_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_7_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_8_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_8_Re <= io_in_8_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_8_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_8_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_8_Im <= io_in_8_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_8_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_9_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_9_Re <= io_in_9_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_9_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_9_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_9_Im <= io_in_9_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_9_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_10_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_10_Re <= io_in_10_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_10_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_10_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_10_Im <= io_in_10_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_10_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_11_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_11_Re <= io_in_11_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_11_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_11_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_11_Im <= io_in_11_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_11_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_12_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_12_Re <= io_in_12_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_12_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_12_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_12_Im <= io_in_12_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_12_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_13_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_13_Re <= io_in_13_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_13_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_13_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_13_Im <= io_in_13_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_13_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_14_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_14_Re <= io_in_14_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_14_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_14_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_14_Im <= io_in_14_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_14_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_15_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_15_Re <= io_in_15_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_15_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_15_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_15_Im <= io_in_15_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_15_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_16_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_16_Re <= io_in_16_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_16_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_16_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_16_Im <= io_in_16_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_16_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_17_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_17_Re <= io_in_17_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_17_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_17_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_17_Im <= io_in_17_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_17_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_18_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_18_Re <= io_in_18_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_18_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_18_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_18_Im <= io_in_18_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_18_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_19_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_19_Re <= io_in_19_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_19_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_19_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_19_Im <= io_in_19_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_19_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_20_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_20_Re <= io_in_20_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_20_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_20_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_20_Im <= io_in_20_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_20_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_21_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_21_Re <= io_in_21_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_21_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_21_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_21_Im <= io_in_21_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_21_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_22_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_22_Re <= io_in_22_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_22_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_22_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_22_Im <= io_in_22_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_22_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_23_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_23_Re <= io_in_23_Re; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_23_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_0_23_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_0_23_Im <= io_in_23_Im; // @[FFTDesigns.scala 2969:38]
    end else begin
      input_delay_registers_0_23_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_0_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_0_Re <= input_delay_registers_0_0_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_0_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_0_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_0_Im <= input_delay_registers_0_0_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_0_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_1_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_1_Re <= input_delay_registers_0_1_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_1_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_1_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_1_Im <= input_delay_registers_0_1_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_1_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_2_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_2_Re <= input_delay_registers_0_2_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_2_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_2_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_2_Im <= input_delay_registers_0_2_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_2_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_3_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_3_Re <= input_delay_registers_0_3_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_3_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_3_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_3_Im <= input_delay_registers_0_3_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_3_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_4_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_4_Re <= input_delay_registers_0_4_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_4_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_4_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_4_Im <= input_delay_registers_0_4_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_4_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_5_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_5_Re <= input_delay_registers_0_5_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_5_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_5_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_5_Im <= input_delay_registers_0_5_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_5_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_6_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_6_Re <= input_delay_registers_0_6_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_6_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_6_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_6_Im <= input_delay_registers_0_6_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_6_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_7_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_7_Re <= input_delay_registers_0_7_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_7_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_7_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_7_Im <= input_delay_registers_0_7_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_7_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_8_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_8_Re <= input_delay_registers_0_8_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_8_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_8_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_8_Im <= input_delay_registers_0_8_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_8_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_9_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_9_Re <= input_delay_registers_0_9_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_9_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_9_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_9_Im <= input_delay_registers_0_9_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_9_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_10_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_10_Re <= input_delay_registers_0_10_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_10_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_10_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_10_Im <= input_delay_registers_0_10_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_10_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_11_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_11_Re <= input_delay_registers_0_11_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_11_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_11_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_11_Im <= input_delay_registers_0_11_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_11_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_12_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_12_Re <= input_delay_registers_0_12_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_12_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_12_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_12_Im <= input_delay_registers_0_12_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_12_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_13_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_13_Re <= input_delay_registers_0_13_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_13_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_13_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_13_Im <= input_delay_registers_0_13_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_13_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_14_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_14_Re <= input_delay_registers_0_14_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_14_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_14_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_14_Im <= input_delay_registers_0_14_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_14_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_15_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_15_Re <= input_delay_registers_0_15_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_15_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_15_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_15_Im <= input_delay_registers_0_15_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_15_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_16_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_16_Re <= input_delay_registers_0_16_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_16_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_16_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_16_Im <= input_delay_registers_0_16_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_16_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_17_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_17_Re <= input_delay_registers_0_17_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_17_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_17_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_17_Im <= input_delay_registers_0_17_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_17_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_18_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_18_Re <= input_delay_registers_0_18_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_18_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_18_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_18_Im <= input_delay_registers_0_18_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_18_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_19_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_19_Re <= input_delay_registers_0_19_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_19_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_19_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_19_Im <= input_delay_registers_0_19_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_19_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_20_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_20_Re <= input_delay_registers_0_20_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_20_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_20_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_20_Im <= input_delay_registers_0_20_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_20_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_21_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_21_Re <= input_delay_registers_0_21_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_21_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_21_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_21_Im <= input_delay_registers_0_21_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_21_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_22_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_22_Re <= input_delay_registers_0_22_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_22_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_22_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_22_Im <= input_delay_registers_0_22_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_22_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_23_Re <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_23_Re <= input_delay_registers_0_23_Re; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_23_Re <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2834:42]
      input_delay_registers_1_23_Im <= 32'h0; // @[FFTDesigns.scala 2834:42]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      input_delay_registers_1_23_Im <= input_delay_registers_0_23_Im; // @[FFTDesigns.scala 2971:38]
    end else begin
      input_delay_registers_1_23_Im <= 32'h0; // @[FFTDesigns.scala 2996:31]
    end
    if (reset) begin // @[FFTDesigns.scala 2912:25]
      cnt2 <= 3'h0; // @[FFTDesigns.scala 2912:25]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      if (cnt2 == 3'h5 & cnt == 2'h3) begin // @[FFTDesigns.scala 2922:69]
        cnt2 <= 3'h0; // @[FFTDesigns.scala 2923:16]
      end else if (_T_3) begin // @[FFTDesigns.scala 2926:47]
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2928:16]
      end else begin
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2931:16]
      end
    end else begin
      cnt2 <= 3'h0; // @[FFTDesigns.scala 3019:14]
    end
    if (reset) begin // @[FFTDesigns.scala 2913:24]
      cnt <= 2'h0; // @[FFTDesigns.scala 2913:24]
    end else if (M0_0_re) begin // @[FFTDesigns.scala 2914:33]
      if (cnt2 == 3'h5 & cnt == 2'h3) begin // @[FFTDesigns.scala 2922:69]
        cnt <= 2'h0; // @[FFTDesigns.scala 2924:15]
      end else if (!(_T_3)) begin // @[FFTDesigns.scala 2926:47]
        cnt <= _GEN_0;
      end
    end else begin
      cnt <= 2'h0; // @[FFTDesigns.scala 3018:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  input_delay_registers_0_0_Re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  input_delay_registers_0_0_Im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  input_delay_registers_0_1_Re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  input_delay_registers_0_1_Im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  input_delay_registers_0_2_Re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  input_delay_registers_0_2_Im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  input_delay_registers_0_3_Re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  input_delay_registers_0_3_Im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  input_delay_registers_0_4_Re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  input_delay_registers_0_4_Im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  input_delay_registers_0_5_Re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  input_delay_registers_0_5_Im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  input_delay_registers_0_6_Re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  input_delay_registers_0_6_Im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  input_delay_registers_0_7_Re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  input_delay_registers_0_7_Im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  input_delay_registers_0_8_Re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  input_delay_registers_0_8_Im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  input_delay_registers_0_9_Re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  input_delay_registers_0_9_Im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  input_delay_registers_0_10_Re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  input_delay_registers_0_10_Im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  input_delay_registers_0_11_Re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  input_delay_registers_0_11_Im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  input_delay_registers_0_12_Re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  input_delay_registers_0_12_Im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  input_delay_registers_0_13_Re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  input_delay_registers_0_13_Im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  input_delay_registers_0_14_Re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  input_delay_registers_0_14_Im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  input_delay_registers_0_15_Re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  input_delay_registers_0_15_Im = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  input_delay_registers_0_16_Re = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  input_delay_registers_0_16_Im = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  input_delay_registers_0_17_Re = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  input_delay_registers_0_17_Im = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  input_delay_registers_0_18_Re = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  input_delay_registers_0_18_Im = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  input_delay_registers_0_19_Re = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  input_delay_registers_0_19_Im = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  input_delay_registers_0_20_Re = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  input_delay_registers_0_20_Im = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  input_delay_registers_0_21_Re = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  input_delay_registers_0_21_Im = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  input_delay_registers_0_22_Re = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  input_delay_registers_0_22_Im = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  input_delay_registers_0_23_Re = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  input_delay_registers_0_23_Im = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  input_delay_registers_1_0_Re = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  input_delay_registers_1_0_Im = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  input_delay_registers_1_1_Re = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  input_delay_registers_1_1_Im = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  input_delay_registers_1_2_Re = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  input_delay_registers_1_2_Im = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  input_delay_registers_1_3_Re = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  input_delay_registers_1_3_Im = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  input_delay_registers_1_4_Re = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  input_delay_registers_1_4_Im = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  input_delay_registers_1_5_Re = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  input_delay_registers_1_5_Im = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  input_delay_registers_1_6_Re = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  input_delay_registers_1_6_Im = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  input_delay_registers_1_7_Re = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  input_delay_registers_1_7_Im = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  input_delay_registers_1_8_Re = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  input_delay_registers_1_8_Im = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  input_delay_registers_1_9_Re = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  input_delay_registers_1_9_Im = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  input_delay_registers_1_10_Re = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  input_delay_registers_1_10_Im = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  input_delay_registers_1_11_Re = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  input_delay_registers_1_11_Im = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  input_delay_registers_1_12_Re = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  input_delay_registers_1_12_Im = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  input_delay_registers_1_13_Re = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  input_delay_registers_1_13_Im = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  input_delay_registers_1_14_Re = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  input_delay_registers_1_14_Im = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  input_delay_registers_1_15_Re = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  input_delay_registers_1_15_Im = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  input_delay_registers_1_16_Re = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  input_delay_registers_1_16_Im = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  input_delay_registers_1_17_Re = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  input_delay_registers_1_17_Im = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  input_delay_registers_1_18_Re = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  input_delay_registers_1_18_Im = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  input_delay_registers_1_19_Re = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  input_delay_registers_1_19_Im = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  input_delay_registers_1_20_Re = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  input_delay_registers_1_20_Im = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  input_delay_registers_1_21_Re = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  input_delay_registers_1_21_Im = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  input_delay_registers_1_22_Re = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  input_delay_registers_1_22_Im = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  input_delay_registers_1_23_Re = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  input_delay_registers_1_23_Im = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  cnt2 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  cnt = _RAND_98[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TwiddleFactorROM_mr(
  input  [6:0]  io_in_addr,
  output [31:0] io_out_data_1_Re,
  output [31:0] io_out_data_1_Im,
  output [31:0] io_out_data_2_Re,
  output [31:0] io_out_data_2_Im,
  output [31:0] io_out_data_4_Re,
  output [31:0] io_out_data_4_Im,
  output [31:0] io_out_data_5_Re,
  output [31:0] io_out_data_5_Im,
  output [31:0] io_out_data_7_Re,
  output [31:0] io_out_data_7_Im,
  output [31:0] io_out_data_8_Re,
  output [31:0] io_out_data_8_Im,
  output [31:0] io_out_data_10_Re,
  output [31:0] io_out_data_10_Im,
  output [31:0] io_out_data_11_Re,
  output [31:0] io_out_data_11_Im,
  output [31:0] io_out_data_13_Re,
  output [31:0] io_out_data_13_Im,
  output [31:0] io_out_data_14_Re,
  output [31:0] io_out_data_14_Im,
  output [31:0] io_out_data_16_Re,
  output [31:0] io_out_data_16_Im,
  output [31:0] io_out_data_17_Re,
  output [31:0] io_out_data_17_Im,
  output [31:0] io_out_data_19_Re,
  output [31:0] io_out_data_19_Im,
  output [31:0] io_out_data_20_Re,
  output [31:0] io_out_data_20_Im,
  output [31:0] io_out_data_22_Re,
  output [31:0] io_out_data_22_Im,
  output [31:0] io_out_data_23_Re,
  output [31:0] io_out_data_23_Im
);
  wire [31:0] _GEN_9 = 2'h1 == io_in_addr[1:0] ? 32'h3f5db3d6 : 32'h3f800000; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_10 = 2'h2 == io_in_addr[1:0] ? 32'h3f000000 : _GEN_9; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_13 = 2'h1 == io_in_addr[1:0] ? 32'hbefffffc : 32'h80800000; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_14 = 2'h2 == io_in_addr[1:0] ? 32'hbf5db3d6 : _GEN_13; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_17 = 2'h1 == io_in_addr[1:0] ? 32'h3f000000 : 32'h3f800000; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_18 = 2'h2 == io_in_addr[1:0] ? 32'hbefffffc : _GEN_17; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_21 = 2'h1 == io_in_addr[1:0] ? 32'hbf5db3d6 : 32'h80800000; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_22 = 2'h2 == io_in_addr[1:0] ? 32'hbf5db3d6 : _GEN_21; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_33 = 2'h1 == io_in_addr[1:0] ? 32'h3f54db30 : 32'h3f7f73ae; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_34 = 2'h2 == io_in_addr[1:0] ? 32'h3ee273a8 : _GEN_33; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_37 = 2'h1 == io_in_addr[1:0] ? 32'hbf0e39d8 : 32'hbd85f210; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_38 = 2'h2 == io_in_addr[1:0] ? 32'hbf659972 : _GEN_37; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_41 = 2'h1 == io_in_addr[1:0] ? 32'h3ec3ef14 : 32'h3f7dcf54; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_42 = 2'h2 == io_in_addr[1:0] ? 32'hbf1bd7c8 : _GEN_41; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_45 = 2'h1 == io_in_addr[1:0] ? 32'hbf6c835e : 32'hbe05a8a8; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_46 = 2'h2 == io_in_addr[1:0] ? 32'hbf4b1934 : _GEN_45; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_57 = 2'h1 == io_in_addr[1:0] ? 32'h3f4b1934 : 32'h3f7dcf54; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_58 = 2'h2 == io_in_addr[1:0] ? 32'h3ec3ef14 : _GEN_57; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_61 = 2'h1 == io_in_addr[1:0] ? 32'hbf1bd7c8 : 32'hbe05a8a8; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_62 = 2'h2 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_61; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_65 = 2'h1 == io_in_addr[1:0] ? 32'h3e8483ec : 32'h3f7746ea; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_66 = 2'h2 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_65; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_69 = 2'h1 == io_in_addr[1:0] ? 32'hbf7746ea : 32'hbe8483ec; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_70 = 2'h2 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_69; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_81 = 2'h1 == io_in_addr[1:0] ? 32'h3f407892 : 32'h3f7b14be; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_82 = 2'h2 == io_in_addr[1:0] ? 32'h3ea493b4 : _GEN_81; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_85 = 2'h1 == io_in_addr[1:0] ? 32'hbf28cae2 : 32'hbe47c5c0; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_86 = 2'h2 == io_in_addr[1:0] ? 32'hbf726a02 : _GEN_85; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_89 = 2'h1 == io_in_addr[1:0] ? 32'h3e05a8a8 : 32'h3f6c835e; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_90 = 2'h2 == io_in_addr[1:0] ? 32'hbf4b1934 : _GEN_89; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_93 = 2'h1 == io_in_addr[1:0] ? 32'hbf7dcf54 : 32'hbec3ef14; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_94 = 2'h2 == io_in_addr[1:0] ? 32'hbf1bd7c8 : _GEN_93; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_105 = 2'h1 == io_in_addr[1:0] ? 32'h3f3504f2 : 32'h3f7746ea; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_106 = 2'h2 == io_in_addr[1:0] ? 32'h3e8483ec : _GEN_105; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_109 = 2'h1 == io_in_addr[1:0] ? 32'hbf3504f2 : 32'hbe8483ec; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_110 = 2'h2 == io_in_addr[1:0] ? 32'hbf7746ea : _GEN_109; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_113 = 2'h1 == io_in_addr[1:0] ? 32'h248d3131 : 32'h3f5db3d6; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_114 = 2'h2 == io_in_addr[1:0] ? 32'hbf5db3d6 : _GEN_113; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_117 = 2'h1 == io_in_addr[1:0] ? 32'hbf800000 : 32'hbefffffc; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_118 = 2'h2 == io_in_addr[1:0] ? 32'hbf000000 : _GEN_117; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_129 = 2'h1 == io_in_addr[1:0] ? 32'h3f28cae2 : 32'h3f726a02; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_130 = 2'h2 == io_in_addr[1:0] ? 32'h3e47c5c0 : _GEN_129; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_133 = 2'h1 == io_in_addr[1:0] ? 32'hbf407892 : 32'hbea493b4; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_134 = 2'h2 == io_in_addr[1:0] ? 32'hbf7b14be : _GEN_133; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_137 = 2'h1 == io_in_addr[1:0] ? 32'hbe05a8a8 : 32'h3f4b1934; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_138 = 2'h2 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_137; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_141 = 2'h1 == io_in_addr[1:0] ? 32'hbf7dcf54 : 32'hbf1bd7c8; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_142 = 2'h2 == io_in_addr[1:0] ? 32'hbec3ef14 : _GEN_141; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_153 = 2'h1 == io_in_addr[1:0] ? 32'h3f1bd7c8 : 32'h3f6c835e; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_154 = 2'h2 == io_in_addr[1:0] ? 32'h3e05a8a8 : _GEN_153; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_157 = 2'h1 == io_in_addr[1:0] ? 32'hbf4b1934 : 32'hbec3ef14; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_158 = 2'h2 == io_in_addr[1:0] ? 32'hbf7dcf54 : _GEN_157; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_161 = 2'h1 == io_in_addr[1:0] ? 32'hbe8483ec : 32'h3f3504f2; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_162 = 2'h2 == io_in_addr[1:0] ? 32'hbf7746ea : _GEN_161; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_165 = 2'h1 == io_in_addr[1:0] ? 32'hbf7746ea : 32'hbf3504f2; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_166 = 2'h2 == io_in_addr[1:0] ? 32'hbe8483ec : _GEN_165; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_177 = 2'h1 == io_in_addr[1:0] ? 32'h3f0e39d8 : 32'h3f659972; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_178 = 2'h2 == io_in_addr[1:0] ? 32'h3d85f210 : _GEN_177; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_181 = 2'h1 == io_in_addr[1:0] ? 32'hbf54db30 : 32'hbee273a8; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_182 = 2'h2 == io_in_addr[1:0] ? 32'hbf7f73ae : _GEN_181; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_185 = 2'h1 == io_in_addr[1:0] ? 32'hbec3ef14 : 32'h3f1bd7c8; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_186 = 2'h2 == io_in_addr[1:0] ? 32'hbf7dcf54 : _GEN_185; // @[FFTDesigns.scala 2084:{25,25}]
  wire [31:0] _GEN_189 = 2'h1 == io_in_addr[1:0] ? 32'hbf6c835e : 32'hbf4b1934; // @[FFTDesigns.scala 2085:{25,25}]
  wire [31:0] _GEN_190 = 2'h2 == io_in_addr[1:0] ? 32'hbe05a8a8 : _GEN_189; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_1_Re = 2'h3 == io_in_addr[1:0] ? 32'h248d3131 : _GEN_10; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_1_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_14; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_2_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf800000 : _GEN_18; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_2_Im = 2'h3 == io_in_addr[1:0] ? 32'ha50d3131 : _GEN_22; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_4_Re = 2'h3 == io_in_addr[1:0] ? 32'hbd85f210 : _GEN_34; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_4_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf7f73ae : _GEN_38; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_5_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf7dcf54 : _GEN_42; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_5_Im = 2'h3 == io_in_addr[1:0] ? 32'h3e05a8a8 : _GEN_46; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_7_Re = 2'h3 == io_in_addr[1:0] ? 32'hbe05a8a8 : _GEN_58; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_7_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf7dcf54 : _GEN_62; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_8_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf7746ea : _GEN_66; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_8_Im = 2'h3 == io_in_addr[1:0] ? 32'h3e8483ec : _GEN_70; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_10_Re = 2'h3 == io_in_addr[1:0] ? 32'hbe47c5c0 : _GEN_82; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_10_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf7b14be : _GEN_86; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_11_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_90; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_11_Im = 2'h3 == io_in_addr[1:0] ? 32'h3ec3ef14 : _GEN_94; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_13_Re = 2'h3 == io_in_addr[1:0] ? 32'hbe8483ec : _GEN_106; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_13_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf7746ea : _GEN_110; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_14_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf5db3d6 : _GEN_114; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_14_Im = 2'h3 == io_in_addr[1:0] ? 32'h3efffffc : _GEN_118; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_16_Re = 2'h3 == io_in_addr[1:0] ? 32'hbea493b4 : _GEN_130; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_16_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf726a02 : _GEN_134; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_17_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf4b1934 : _GEN_138; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_17_Im = 2'h3 == io_in_addr[1:0] ? 32'h3f1bd7c8 : _GEN_142; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_19_Re = 2'h3 == io_in_addr[1:0] ? 32'hbec3ef14 : _GEN_154; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_19_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf6c835e : _GEN_158; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_20_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf3504f2 : _GEN_162; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_20_Im = 2'h3 == io_in_addr[1:0] ? 32'h3f3504f2 : _GEN_166; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_22_Re = 2'h3 == io_in_addr[1:0] ? 32'hbee273a8 : _GEN_178; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_22_Im = 2'h3 == io_in_addr[1:0] ? 32'hbf659972 : _GEN_182; // @[FFTDesigns.scala 2085:{25,25}]
  assign io_out_data_23_Re = 2'h3 == io_in_addr[1:0] ? 32'hbf1bd7c8 : _GEN_186; // @[FFTDesigns.scala 2084:{25,25}]
  assign io_out_data_23_Im = 2'h3 == io_in_addr[1:0] ? 32'h3f4b1934 : _GEN_190; // @[FFTDesigns.scala 2085:{25,25}]
endmodule
module TwiddleFactorsStreamed_mr_v2(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input  [31:0] io_in_16_Re,
  input  [31:0] io_in_16_Im,
  input  [31:0] io_in_17_Re,
  input  [31:0] io_in_17_Im,
  input  [31:0] io_in_18_Re,
  input  [31:0] io_in_18_Im,
  input  [31:0] io_in_19_Re,
  input  [31:0] io_in_19_Im,
  input  [31:0] io_in_20_Re,
  input  [31:0] io_in_20_Im,
  input  [31:0] io_in_21_Re,
  input  [31:0] io_in_21_Im,
  input  [31:0] io_in_22_Re,
  input  [31:0] io_in_22_Im,
  input  [31:0] io_in_23_Re,
  input  [31:0] io_in_23_Im,
  input         io_in_en_0,
  input         io_in_en_1,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im,
  output [31:0] io_out_16_Re,
  output [31:0] io_out_16_Im,
  output [31:0] io_out_17_Re,
  output [31:0] io_out_17_Im,
  output [31:0] io_out_18_Re,
  output [31:0] io_out_18_Im,
  output [31:0] io_out_19_Re,
  output [31:0] io_out_19_Im,
  output [31:0] io_out_20_Re,
  output [31:0] io_out_20_Im,
  output [31:0] io_out_21_Re,
  output [31:0] io_out_21_Im,
  output [31:0] io_out_22_Re,
  output [31:0] io_out_22_Im,
  output [31:0] io_out_23_Re,
  output [31:0] io_out_23_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] TwiddleFactorROM_mr_io_in_addr; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_1_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_1_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_2_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_2_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_4_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_4_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_5_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_5_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_7_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_7_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_8_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_8_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_10_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_10_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_11_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_11_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_13_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_13_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_14_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_14_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_16_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_16_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_17_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_17_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_19_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_19_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_20_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_20_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_22_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_22_Im; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_23_Re; // @[FFTDesigns.scala 2314:26]
  wire [31:0] TwiddleFactorROM_mr_io_out_data_23_Im; // @[FFTDesigns.scala 2314:26]
  wire  FPComplexMult_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_1_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_1_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_2_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_2_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_3_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_3_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_4_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_4_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_5_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_5_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_6_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_6_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_7_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_7_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_8_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_8_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_9_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_9_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_10_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_10_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_11_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_11_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_12_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_12_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_12_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_12_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_12_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_12_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_13_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_13_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_13_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_13_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_13_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_13_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_14_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_14_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_14_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_14_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_14_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_14_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_15_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_15_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_15_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_15_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_15_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_15_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_16_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_16_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_16_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_16_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_16_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_16_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_16_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_16_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_17_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_17_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_17_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_17_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_17_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_17_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_17_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_17_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_18_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_18_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_18_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_18_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_18_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_18_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_18_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_18_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_19_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_19_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_19_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_19_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_19_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_19_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_19_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_19_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_20_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_20_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_20_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_20_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_20_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_20_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_20_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_20_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_21_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_21_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_21_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_21_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_21_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_21_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_21_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_21_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_22_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_22_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_22_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_22_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_22_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_22_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_22_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_22_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_23_clock; // @[FFTDesigns.scala 2330:30]
  wire  FPComplexMult_23_reset; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_23_io_in_a_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_23_io_in_a_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_23_io_in_b_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_23_io_in_b_Im; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_23_io_out_s_Re; // @[FFTDesigns.scala 2330:30]
  wire [31:0] FPComplexMult_23_io_out_s_Im; // @[FFTDesigns.scala 2330:30]
  reg [1:0] cnt; // @[FFTDesigns.scala 2322:24]
  reg [2:0] cnt2; // @[FFTDesigns.scala 2323:25]
  wire [1:0] _T = {io_in_en_1,io_in_en_0}; // @[FFTDesigns.scala 2324:21]
  wire  _T_1 = |_T; // @[FFTDesigns.scala 2324:28]
  wire [2:0] _cnt2_T_1 = cnt2 + 3'h1; // @[FFTDesigns.scala 2339:24]
  wire [1:0] _cnt_T_1 = cnt + 2'h1; // @[FFTDesigns.scala 2341:22]
  TwiddleFactorROM_mr TwiddleFactorROM_mr ( // @[FFTDesigns.scala 2314:26]
    .io_in_addr(TwiddleFactorROM_mr_io_in_addr),
    .io_out_data_1_Re(TwiddleFactorROM_mr_io_out_data_1_Re),
    .io_out_data_1_Im(TwiddleFactorROM_mr_io_out_data_1_Im),
    .io_out_data_2_Re(TwiddleFactorROM_mr_io_out_data_2_Re),
    .io_out_data_2_Im(TwiddleFactorROM_mr_io_out_data_2_Im),
    .io_out_data_4_Re(TwiddleFactorROM_mr_io_out_data_4_Re),
    .io_out_data_4_Im(TwiddleFactorROM_mr_io_out_data_4_Im),
    .io_out_data_5_Re(TwiddleFactorROM_mr_io_out_data_5_Re),
    .io_out_data_5_Im(TwiddleFactorROM_mr_io_out_data_5_Im),
    .io_out_data_7_Re(TwiddleFactorROM_mr_io_out_data_7_Re),
    .io_out_data_7_Im(TwiddleFactorROM_mr_io_out_data_7_Im),
    .io_out_data_8_Re(TwiddleFactorROM_mr_io_out_data_8_Re),
    .io_out_data_8_Im(TwiddleFactorROM_mr_io_out_data_8_Im),
    .io_out_data_10_Re(TwiddleFactorROM_mr_io_out_data_10_Re),
    .io_out_data_10_Im(TwiddleFactorROM_mr_io_out_data_10_Im),
    .io_out_data_11_Re(TwiddleFactorROM_mr_io_out_data_11_Re),
    .io_out_data_11_Im(TwiddleFactorROM_mr_io_out_data_11_Im),
    .io_out_data_13_Re(TwiddleFactorROM_mr_io_out_data_13_Re),
    .io_out_data_13_Im(TwiddleFactorROM_mr_io_out_data_13_Im),
    .io_out_data_14_Re(TwiddleFactorROM_mr_io_out_data_14_Re),
    .io_out_data_14_Im(TwiddleFactorROM_mr_io_out_data_14_Im),
    .io_out_data_16_Re(TwiddleFactorROM_mr_io_out_data_16_Re),
    .io_out_data_16_Im(TwiddleFactorROM_mr_io_out_data_16_Im),
    .io_out_data_17_Re(TwiddleFactorROM_mr_io_out_data_17_Re),
    .io_out_data_17_Im(TwiddleFactorROM_mr_io_out_data_17_Im),
    .io_out_data_19_Re(TwiddleFactorROM_mr_io_out_data_19_Re),
    .io_out_data_19_Im(TwiddleFactorROM_mr_io_out_data_19_Im),
    .io_out_data_20_Re(TwiddleFactorROM_mr_io_out_data_20_Re),
    .io_out_data_20_Im(TwiddleFactorROM_mr_io_out_data_20_Im),
    .io_out_data_22_Re(TwiddleFactorROM_mr_io_out_data_22_Re),
    .io_out_data_22_Im(TwiddleFactorROM_mr_io_out_data_22_Im),
    .io_out_data_23_Re(TwiddleFactorROM_mr_io_out_data_23_Re),
    .io_out_data_23_Im(TwiddleFactorROM_mr_io_out_data_23_Im)
  );
  FPComplexMult FPComplexMult ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_clock),
    .reset(FPComplexMult_reset),
    .io_in_a_Re(FPComplexMult_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_1 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_1_clock),
    .reset(FPComplexMult_1_reset),
    .io_in_a_Re(FPComplexMult_1_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_1_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_1_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_1_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_1_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_1_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_2 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_2_clock),
    .reset(FPComplexMult_2_reset),
    .io_in_a_Re(FPComplexMult_2_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_2_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_2_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_2_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_2_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_2_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_3 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_3_clock),
    .reset(FPComplexMult_3_reset),
    .io_in_a_Re(FPComplexMult_3_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_3_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_3_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_3_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_3_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_3_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_4 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_4_clock),
    .reset(FPComplexMult_4_reset),
    .io_in_a_Re(FPComplexMult_4_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_4_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_4_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_4_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_4_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_4_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_5 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_5_clock),
    .reset(FPComplexMult_5_reset),
    .io_in_a_Re(FPComplexMult_5_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_5_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_5_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_5_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_5_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_5_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_6 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_6_clock),
    .reset(FPComplexMult_6_reset),
    .io_in_a_Re(FPComplexMult_6_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_6_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_6_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_6_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_6_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_6_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_7 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_7_clock),
    .reset(FPComplexMult_7_reset),
    .io_in_a_Re(FPComplexMult_7_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_7_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_7_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_7_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_7_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_7_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_8 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_8_clock),
    .reset(FPComplexMult_8_reset),
    .io_in_a_Re(FPComplexMult_8_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_8_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_8_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_8_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_8_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_8_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_9 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_9_clock),
    .reset(FPComplexMult_9_reset),
    .io_in_a_Re(FPComplexMult_9_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_9_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_9_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_9_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_9_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_9_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_10 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_10_clock),
    .reset(FPComplexMult_10_reset),
    .io_in_a_Re(FPComplexMult_10_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_10_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_10_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_10_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_10_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_10_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_11 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_11_clock),
    .reset(FPComplexMult_11_reset),
    .io_in_a_Re(FPComplexMult_11_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_11_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_11_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_11_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_11_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_11_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_12 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_12_clock),
    .reset(FPComplexMult_12_reset),
    .io_in_a_Re(FPComplexMult_12_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_12_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_12_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_12_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_12_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_12_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_13 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_13_clock),
    .reset(FPComplexMult_13_reset),
    .io_in_a_Re(FPComplexMult_13_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_13_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_13_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_13_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_13_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_13_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_14 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_14_clock),
    .reset(FPComplexMult_14_reset),
    .io_in_a_Re(FPComplexMult_14_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_14_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_14_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_14_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_14_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_14_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_15 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_15_clock),
    .reset(FPComplexMult_15_reset),
    .io_in_a_Re(FPComplexMult_15_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_15_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_15_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_15_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_15_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_15_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_16 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_16_clock),
    .reset(FPComplexMult_16_reset),
    .io_in_a_Re(FPComplexMult_16_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_16_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_16_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_16_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_16_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_16_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_17 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_17_clock),
    .reset(FPComplexMult_17_reset),
    .io_in_a_Re(FPComplexMult_17_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_17_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_17_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_17_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_17_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_17_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_18 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_18_clock),
    .reset(FPComplexMult_18_reset),
    .io_in_a_Re(FPComplexMult_18_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_18_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_18_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_18_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_18_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_18_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_19 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_19_clock),
    .reset(FPComplexMult_19_reset),
    .io_in_a_Re(FPComplexMult_19_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_19_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_19_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_19_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_19_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_19_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_20 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_20_clock),
    .reset(FPComplexMult_20_reset),
    .io_in_a_Re(FPComplexMult_20_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_20_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_20_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_20_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_20_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_20_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_21 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_21_clock),
    .reset(FPComplexMult_21_reset),
    .io_in_a_Re(FPComplexMult_21_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_21_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_21_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_21_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_21_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_21_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_22 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_22_clock),
    .reset(FPComplexMult_22_reset),
    .io_in_a_Re(FPComplexMult_22_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_22_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_22_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_22_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_22_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_22_io_out_s_Im)
  );
  FPComplexMult FPComplexMult_23 ( // @[FFTDesigns.scala 2330:30]
    .clock(FPComplexMult_23_clock),
    .reset(FPComplexMult_23_reset),
    .io_in_a_Re(FPComplexMult_23_io_in_a_Re),
    .io_in_a_Im(FPComplexMult_23_io_in_a_Im),
    .io_in_b_Re(FPComplexMult_23_io_in_b_Re),
    .io_in_b_Im(FPComplexMult_23_io_in_b_Im),
    .io_out_s_Re(FPComplexMult_23_io_out_s_Re),
    .io_out_s_Im(FPComplexMult_23_io_out_s_Im)
  );
  assign io_out_0_Re = FPComplexMult_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_0_Im = FPComplexMult_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_1_Re = FPComplexMult_1_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_1_Im = FPComplexMult_1_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_2_Re = FPComplexMult_2_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_2_Im = FPComplexMult_2_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_3_Re = FPComplexMult_3_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_3_Im = FPComplexMult_3_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_4_Re = FPComplexMult_4_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_4_Im = FPComplexMult_4_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_5_Re = FPComplexMult_5_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_5_Im = FPComplexMult_5_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_6_Re = FPComplexMult_6_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_6_Im = FPComplexMult_6_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_7_Re = FPComplexMult_7_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_7_Im = FPComplexMult_7_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_8_Re = FPComplexMult_8_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_8_Im = FPComplexMult_8_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_9_Re = FPComplexMult_9_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_9_Im = FPComplexMult_9_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_10_Re = FPComplexMult_10_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_10_Im = FPComplexMult_10_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_11_Re = FPComplexMult_11_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_11_Im = FPComplexMult_11_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_12_Re = FPComplexMult_12_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_12_Im = FPComplexMult_12_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_13_Re = FPComplexMult_13_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_13_Im = FPComplexMult_13_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_14_Re = FPComplexMult_14_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_14_Im = FPComplexMult_14_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_15_Re = FPComplexMult_15_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_15_Im = FPComplexMult_15_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_16_Re = FPComplexMult_16_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_16_Im = FPComplexMult_16_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_17_Re = FPComplexMult_17_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_17_Im = FPComplexMult_17_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_18_Re = FPComplexMult_18_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_18_Im = FPComplexMult_18_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_19_Re = FPComplexMult_19_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_19_Im = FPComplexMult_19_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_20_Re = FPComplexMult_20_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_20_Im = FPComplexMult_20_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_21_Re = FPComplexMult_21_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_21_Im = FPComplexMult_21_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_22_Re = FPComplexMult_22_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_22_Im = FPComplexMult_22_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign io_out_23_Re = FPComplexMult_23_io_out_s_Re; // @[FFTDesigns.scala 2357:19]
  assign io_out_23_Im = FPComplexMult_23_io_out_s_Im; // @[FFTDesigns.scala 2357:19]
  assign TwiddleFactorROM_mr_io_in_addr = {{5'd0}, cnt}; // @[FFTDesigns.scala 2359:24]
  assign FPComplexMult_clock = clock;
  assign FPComplexMult_reset = reset;
  assign FPComplexMult_io_in_a_Re = _T_1 ? io_in_0_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_io_in_a_Im = _T_1 ? io_in_0_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_1_clock = clock;
  assign FPComplexMult_1_reset = reset;
  assign FPComplexMult_1_io_in_a_Re = _T_1 ? io_in_1_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_1_io_in_a_Im = _T_1 ? io_in_1_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_1_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_1_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_1_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_1_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_2_clock = clock;
  assign FPComplexMult_2_reset = reset;
  assign FPComplexMult_2_io_in_a_Re = _T_1 ? io_in_2_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_2_io_in_a_Im = _T_1 ? io_in_2_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_2_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_2_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_2_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_2_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_3_clock = clock;
  assign FPComplexMult_3_reset = reset;
  assign FPComplexMult_3_io_in_a_Re = _T_1 ? io_in_3_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_3_io_in_a_Im = _T_1 ? io_in_3_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_3_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_3_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_4_clock = clock;
  assign FPComplexMult_4_reset = reset;
  assign FPComplexMult_4_io_in_a_Re = _T_1 ? io_in_4_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_4_io_in_a_Im = _T_1 ? io_in_4_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_4_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_4_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_4_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_4_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_5_clock = clock;
  assign FPComplexMult_5_reset = reset;
  assign FPComplexMult_5_io_in_a_Re = _T_1 ? io_in_5_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_5_io_in_a_Im = _T_1 ? io_in_5_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_5_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_5_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_5_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_5_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_6_clock = clock;
  assign FPComplexMult_6_reset = reset;
  assign FPComplexMult_6_io_in_a_Re = _T_1 ? io_in_6_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_6_io_in_a_Im = _T_1 ? io_in_6_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_6_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_6_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_7_clock = clock;
  assign FPComplexMult_7_reset = reset;
  assign FPComplexMult_7_io_in_a_Re = _T_1 ? io_in_7_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_7_io_in_a_Im = _T_1 ? io_in_7_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_7_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_7_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_7_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_7_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_8_clock = clock;
  assign FPComplexMult_8_reset = reset;
  assign FPComplexMult_8_io_in_a_Re = _T_1 ? io_in_8_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_8_io_in_a_Im = _T_1 ? io_in_8_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_8_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_8_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_8_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_8_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_9_clock = clock;
  assign FPComplexMult_9_reset = reset;
  assign FPComplexMult_9_io_in_a_Re = _T_1 ? io_in_9_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_9_io_in_a_Im = _T_1 ? io_in_9_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_9_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_9_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_10_clock = clock;
  assign FPComplexMult_10_reset = reset;
  assign FPComplexMult_10_io_in_a_Re = _T_1 ? io_in_10_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_10_io_in_a_Im = _T_1 ? io_in_10_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_10_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_10_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_10_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_10_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_11_clock = clock;
  assign FPComplexMult_11_reset = reset;
  assign FPComplexMult_11_io_in_a_Re = _T_1 ? io_in_11_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_11_io_in_a_Im = _T_1 ? io_in_11_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_11_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_11_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_11_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_11_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_12_clock = clock;
  assign FPComplexMult_12_reset = reset;
  assign FPComplexMult_12_io_in_a_Re = _T_1 ? io_in_12_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_12_io_in_a_Im = _T_1 ? io_in_12_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_12_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_12_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_13_clock = clock;
  assign FPComplexMult_13_reset = reset;
  assign FPComplexMult_13_io_in_a_Re = _T_1 ? io_in_13_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_13_io_in_a_Im = _T_1 ? io_in_13_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_13_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_13_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_13_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_13_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_14_clock = clock;
  assign FPComplexMult_14_reset = reset;
  assign FPComplexMult_14_io_in_a_Re = _T_1 ? io_in_14_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_14_io_in_a_Im = _T_1 ? io_in_14_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_14_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_14_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_14_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_14_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_15_clock = clock;
  assign FPComplexMult_15_reset = reset;
  assign FPComplexMult_15_io_in_a_Re = _T_1 ? io_in_15_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_15_io_in_a_Im = _T_1 ? io_in_15_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_15_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_15_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_16_clock = clock;
  assign FPComplexMult_16_reset = reset;
  assign FPComplexMult_16_io_in_a_Re = _T_1 ? io_in_16_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_16_io_in_a_Im = _T_1 ? io_in_16_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_16_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_16_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_16_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_16_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_17_clock = clock;
  assign FPComplexMult_17_reset = reset;
  assign FPComplexMult_17_io_in_a_Re = _T_1 ? io_in_17_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_17_io_in_a_Im = _T_1 ? io_in_17_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_17_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_17_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_17_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_17_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_18_clock = clock;
  assign FPComplexMult_18_reset = reset;
  assign FPComplexMult_18_io_in_a_Re = _T_1 ? io_in_18_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_18_io_in_a_Im = _T_1 ? io_in_18_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_18_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_18_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_19_clock = clock;
  assign FPComplexMult_19_reset = reset;
  assign FPComplexMult_19_io_in_a_Re = _T_1 ? io_in_19_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_19_io_in_a_Im = _T_1 ? io_in_19_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_19_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_19_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_19_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_19_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_20_clock = clock;
  assign FPComplexMult_20_reset = reset;
  assign FPComplexMult_20_io_in_a_Re = _T_1 ? io_in_20_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_20_io_in_a_Im = _T_1 ? io_in_20_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_20_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_20_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_20_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_20_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_21_clock = clock;
  assign FPComplexMult_21_reset = reset;
  assign FPComplexMult_21_io_in_a_Re = _T_1 ? io_in_21_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_21_io_in_a_Im = _T_1 ? io_in_21_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_21_io_in_b_Re = _T_1 ? 32'h3f800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_21_io_in_b_Im = _T_1 ? 32'h80800000 : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_22_clock = clock;
  assign FPComplexMult_22_reset = reset;
  assign FPComplexMult_22_io_in_a_Re = _T_1 ? io_in_22_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_22_io_in_a_Im = _T_1 ? io_in_22_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_22_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_22_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_22_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_22_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_23_clock = clock;
  assign FPComplexMult_23_reset = reset;
  assign FPComplexMult_23_io_in_a_Re = _T_1 ? io_in_23_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_23_io_in_a_Im = _T_1 ? io_in_23_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2345:31 2350:31]
  assign FPComplexMult_23_io_in_b_Re = _T_1 ? TwiddleFactorROM_mr_io_out_data_23_Re : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  assign FPComplexMult_23_io_in_b_Im = _T_1 ? TwiddleFactorROM_mr_io_out_data_23_Im : 32'h0; // @[FFTDesigns.scala 2333:32 2346:31 2351:31]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 2322:24]
      cnt <= 2'h0; // @[FFTDesigns.scala 2322:24]
    end else if (_T_1) begin // @[FFTDesigns.scala 2333:32]
      if (cnt2 == 3'h5) begin // @[FFTDesigns.scala 2334:37]
        cnt <= 2'h0; // @[FFTDesigns.scala 2336:15]
      end else if (!(cnt == 2'h3 & cnt2 != 3'h5)) begin // @[FFTDesigns.scala 2337:66]
        cnt <= _cnt_T_1; // @[FFTDesigns.scala 2341:15]
      end
    end else begin
      cnt <= 2'h0; // @[FFTDesigns.scala 2353:13]
    end
    if (reset) begin // @[FFTDesigns.scala 2323:25]
      cnt2 <= 3'h0; // @[FFTDesigns.scala 2323:25]
    end else if (_T_1) begin // @[FFTDesigns.scala 2333:32]
      if (cnt2 == 3'h5) begin // @[FFTDesigns.scala 2334:37]
        cnt2 <= 3'h0; // @[FFTDesigns.scala 2335:16]
      end else if (cnt == 2'h3 & cnt2 != 3'h5) begin // @[FFTDesigns.scala 2337:66]
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2339:16]
      end else begin
        cnt2 <= _cnt2_T_1; // @[FFTDesigns.scala 2342:16]
      end
    end else begin
      cnt2 <= 3'h0; // @[FFTDesigns.scala 2354:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cnt2 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module od_fft96_16_24(
  input         clock,
  input         reset,
  input  [31:0] io_in_0_Re,
  input  [31:0] io_in_0_Im,
  input  [31:0] io_in_1_Re,
  input  [31:0] io_in_1_Im,
  input  [31:0] io_in_2_Re,
  input  [31:0] io_in_2_Im,
  input  [31:0] io_in_3_Re,
  input  [31:0] io_in_3_Im,
  input  [31:0] io_in_4_Re,
  input  [31:0] io_in_4_Im,
  input  [31:0] io_in_5_Re,
  input  [31:0] io_in_5_Im,
  input  [31:0] io_in_6_Re,
  input  [31:0] io_in_6_Im,
  input  [31:0] io_in_7_Re,
  input  [31:0] io_in_7_Im,
  input  [31:0] io_in_8_Re,
  input  [31:0] io_in_8_Im,
  input  [31:0] io_in_9_Re,
  input  [31:0] io_in_9_Im,
  input  [31:0] io_in_10_Re,
  input  [31:0] io_in_10_Im,
  input  [31:0] io_in_11_Re,
  input  [31:0] io_in_11_Im,
  input  [31:0] io_in_12_Re,
  input  [31:0] io_in_12_Im,
  input  [31:0] io_in_13_Re,
  input  [31:0] io_in_13_Im,
  input  [31:0] io_in_14_Re,
  input  [31:0] io_in_14_Im,
  input  [31:0] io_in_15_Re,
  input  [31:0] io_in_15_Im,
  input         io_in_ready,
  output        io_out_validate,
  output [31:0] io_out_0_Re,
  output [31:0] io_out_0_Im,
  output [31:0] io_out_1_Re,
  output [31:0] io_out_1_Im,
  output [31:0] io_out_2_Re,
  output [31:0] io_out_2_Im,
  output [31:0] io_out_3_Re,
  output [31:0] io_out_3_Im,
  output [31:0] io_out_4_Re,
  output [31:0] io_out_4_Im,
  output [31:0] io_out_5_Re,
  output [31:0] io_out_5_Im,
  output [31:0] io_out_6_Re,
  output [31:0] io_out_6_Im,
  output [31:0] io_out_7_Re,
  output [31:0] io_out_7_Im,
  output [31:0] io_out_8_Re,
  output [31:0] io_out_8_Im,
  output [31:0] io_out_9_Re,
  output [31:0] io_out_9_Im,
  output [31:0] io_out_10_Re,
  output [31:0] io_out_10_Im,
  output [31:0] io_out_11_Re,
  output [31:0] io_out_11_Im,
  output [31:0] io_out_12_Re,
  output [31:0] io_out_12_Im,
  output [31:0] io_out_13_Re,
  output [31:0] io_out_13_Im,
  output [31:0] io_out_14_Re,
  output [31:0] io_out_14_Im,
  output [31:0] io_out_15_Re,
  output [31:0] io_out_15_Im
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_REG_INIT
  wire  FFT_sr_v2_streaming_nrv_clock; // @[FFTDesigns.scala 6453:32]
  wire  FFT_sr_v2_streaming_nrv_reset; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_0_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_0_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_1_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_1_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_2_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_2_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_3_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_3_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_4_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_4_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_5_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_5_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_6_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_6_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_7_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_7_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_8_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_8_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_9_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_9_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_10_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_10_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_11_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_11_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_12_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_12_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_13_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_13_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_14_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_14_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_15_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_in_15_Im; // @[FFTDesigns.scala 6453:32]
  wire  FFT_sr_v2_streaming_nrv_io_in_ready; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_0_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_0_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_1_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_1_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_2_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_2_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_3_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_3_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_4_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_4_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_5_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_5_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_6_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_6_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_7_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_7_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_8_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_8_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_9_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_9_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_10_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_10_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_11_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_11_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_12_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_12_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_13_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_13_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_14_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_14_Im; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_15_Re; // @[FFTDesigns.scala 6453:32]
  wire [31:0] FFT_sr_v2_streaming_nrv_io_out_15_Im; // @[FFTDesigns.scala 6453:32]
  wire  DFT_r_v2_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_1_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_1_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_1_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_2_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_2_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_2_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_3_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_3_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_3_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_4_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_4_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_4_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_5_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_5_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_5_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_6_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_6_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_6_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_7_clock; // @[FFTDesigns.scala 6457:32]
  wire  DFT_r_v2_7_reset; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_in_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_in_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_in_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_in_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_in_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_in_2_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_out_0_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_out_0_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_out_1_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_out_1_Im; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_out_2_Re; // @[FFTDesigns.scala 6457:32]
  wire [31:0] DFT_r_v2_7_io_out_2_Im; // @[FFTDesigns.scala 6457:32]
  wire  PermutationsWithStreaming_clock; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_reset; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_0_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_0_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_1_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_1_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_2_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_2_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_3_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_3_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_4_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_4_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_5_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_5_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_6_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_6_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_7_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_7_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_8_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_8_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_9_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_9_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_10_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_10_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_11_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_11_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_12_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_12_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_13_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_13_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_14_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_14_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_15_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_in_15_Im; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_0; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_1; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_2; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_3; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_4; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_5; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_6; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_7; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_8; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_9; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_10; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_11; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_io_in_en_12; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_0_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_0_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_1_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_1_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_2_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_2_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_3_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_3_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_4_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_4_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_5_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_5_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_6_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_6_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_7_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_7_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_8_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_8_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_9_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_9_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_10_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_10_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_11_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_11_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_12_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_12_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_13_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_13_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_14_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_14_Im; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_15_Re; // @[FFTDesigns.scala 6468:32]
  wire [31:0] PermutationsWithStreaming_io_out_15_Im; // @[FFTDesigns.scala 6468:32]
  wire  PermutationsWithStreaming_mr_clock; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_reset; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_0_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_0_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_1_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_1_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_2_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_2_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_3_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_3_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_4_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_4_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_5_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_5_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_6_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_6_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_7_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_7_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_8_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_8_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_9_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_9_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_10_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_10_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_11_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_11_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_12_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_12_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_13_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_13_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_14_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_14_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_15_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_in_15_Im; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_0; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_1; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_2; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_3; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_4; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_5; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_6; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_7; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_8; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_9; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_10; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_11; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_io_in_en_12; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_0_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_0_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_1_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_1_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_2_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_2_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_3_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_3_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_4_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_4_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_5_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_5_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_6_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_6_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_7_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_7_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_8_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_8_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_9_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_9_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_10_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_10_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_11_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_11_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_12_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_12_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_13_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_13_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_14_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_14_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_15_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_15_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_16_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_16_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_17_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_17_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_18_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_18_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_19_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_19_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_20_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_20_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_21_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_21_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_22_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_22_Im; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_23_Re; // @[FFTDesigns.scala 6469:32]
  wire [31:0] PermutationsWithStreaming_mr_io_out_23_Im; // @[FFTDesigns.scala 6469:32]
  wire  PermutationsWithStreaming_mr_1_clock; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_reset; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_0_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_0_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_1_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_1_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_2_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_2_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_3_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_3_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_4_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_4_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_5_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_5_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_6_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_6_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_7_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_7_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_8_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_8_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_9_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_9_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_10_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_10_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_11_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_11_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_12_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_12_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_13_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_13_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_14_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_14_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_15_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_15_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_16_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_16_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_17_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_17_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_18_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_18_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_19_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_19_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_20_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_20_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_21_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_21_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_22_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_22_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_23_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_in_23_Im; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_0; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_1; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_2; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_3; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_4; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_5; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_6; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_7; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_8; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_9; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_10; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_11; // @[FFTDesigns.scala 6470:32]
  wire  PermutationsWithStreaming_mr_1_io_in_en_12; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_0_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_0_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_1_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_1_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_2_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_2_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_3_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_3_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_4_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_4_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_5_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_5_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_6_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_6_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_7_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_7_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_8_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_8_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_9_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_9_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_10_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_10_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_11_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_11_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_12_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_12_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_13_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_13_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_14_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_14_Im; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_15_Re; // @[FFTDesigns.scala 6470:32]
  wire [31:0] PermutationsWithStreaming_mr_1_io_out_15_Im; // @[FFTDesigns.scala 6470:32]
  wire  TwiddleFactorsStreamed_mr_v2_clock; // @[FFTDesigns.scala 6471:32]
  wire  TwiddleFactorsStreamed_mr_v2_reset; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_0_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_0_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_1_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_1_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_2_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_2_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_3_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_3_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_4_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_4_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_5_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_5_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_6_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_6_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_7_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_7_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_8_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_8_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_9_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_9_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_10_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_10_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_11_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_11_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_12_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_12_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_13_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_13_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_14_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_14_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_15_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_15_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_16_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_16_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_17_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_17_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_18_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_18_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_19_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_19_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_20_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_20_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_21_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_21_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_22_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_22_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_23_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_in_23_Im; // @[FFTDesigns.scala 6471:32]
  wire  TwiddleFactorsStreamed_mr_v2_io_in_en_0; // @[FFTDesigns.scala 6471:32]
  wire  TwiddleFactorsStreamed_mr_v2_io_in_en_1; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_0_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_0_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_1_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_1_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_2_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_2_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_3_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_3_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_4_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_4_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_5_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_5_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_6_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_6_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_7_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_7_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_8_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_8_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_9_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_9_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_10_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_10_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_11_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_11_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_12_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_12_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_13_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_13_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_14_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_14_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_15_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_15_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_16_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_16_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_17_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_17_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_18_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_18_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_19_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_19_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_20_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_20_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_21_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_21_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_22_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_22_Im; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_23_Re; // @[FFTDesigns.scala 6471:32]
  wire [31:0] TwiddleFactorsStreamed_mr_v2_io_out_23_Im; // @[FFTDesigns.scala 6471:32]
  reg  DFT_regdelays1_0; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_1; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_2; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_3; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_4; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_5; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_6; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_7; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_8; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_9; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_10; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_11; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_12; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_13; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_14; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_15; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_16; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_17; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_18; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_19; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_20; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_21; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_22; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_23; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_24; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_25; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_26; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_27; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_28; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_29; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_30; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_31; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_32; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_33; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_34; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_35; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays1_36; // @[FFTDesigns.scala 6474:35]
  reg  DFT_regdelays2_0; // @[FFTDesigns.scala 6475:35]
  reg  DFT_regdelays2_1; // @[FFTDesigns.scala 6475:35]
  reg  DFT_regdelays2_2; // @[FFTDesigns.scala 6475:35]
  reg  DFT_regdelays2_3; // @[FFTDesigns.scala 6475:35]
  reg  Twid_regdelays_0; // @[FFTDesigns.scala 6476:35]
  reg  Twid_regdelays_1; // @[FFTDesigns.scala 6476:35]
  reg  Perm_regdelays1_0_0; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_1; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_2; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_3; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_4; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_5; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_6; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_7; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_8; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_9; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_10; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_0_11; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_0; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_1; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_2; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_3; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_4; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_5; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_6; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_7; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_8; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_9; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_10; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_1_11; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_0; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_1; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_2; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_3; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_4; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_5; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_6; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_7; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_8; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_9; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_10; // @[FFTDesigns.scala 6477:36]
  reg  Perm_regdelays1_2_11; // @[FFTDesigns.scala 6477:36]
  reg  out_regdelay; // @[FFTDesigns.scala 6478:33]
  reg [31:0] results_0_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_0_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_1_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_1_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_2_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_2_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_3_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_3_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_4_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_4_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_5_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_5_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_6_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_6_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_7_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_7_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_8_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_8_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_9_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_9_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_10_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_10_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_11_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_11_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_12_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_12_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_13_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_13_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_14_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_14_Im; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_15_Re; // @[FFTDesigns.scala 6479:28]
  reg [31:0] results_15_Im; // @[FFTDesigns.scala 6479:28]
  FFT_sr_v2_streaming_nrv FFT_sr_v2_streaming_nrv ( // @[FFTDesigns.scala 6453:32]
    .clock(FFT_sr_v2_streaming_nrv_clock),
    .reset(FFT_sr_v2_streaming_nrv_reset),
    .io_in_0_Re(FFT_sr_v2_streaming_nrv_io_in_0_Re),
    .io_in_0_Im(FFT_sr_v2_streaming_nrv_io_in_0_Im),
    .io_in_1_Re(FFT_sr_v2_streaming_nrv_io_in_1_Re),
    .io_in_1_Im(FFT_sr_v2_streaming_nrv_io_in_1_Im),
    .io_in_2_Re(FFT_sr_v2_streaming_nrv_io_in_2_Re),
    .io_in_2_Im(FFT_sr_v2_streaming_nrv_io_in_2_Im),
    .io_in_3_Re(FFT_sr_v2_streaming_nrv_io_in_3_Re),
    .io_in_3_Im(FFT_sr_v2_streaming_nrv_io_in_3_Im),
    .io_in_4_Re(FFT_sr_v2_streaming_nrv_io_in_4_Re),
    .io_in_4_Im(FFT_sr_v2_streaming_nrv_io_in_4_Im),
    .io_in_5_Re(FFT_sr_v2_streaming_nrv_io_in_5_Re),
    .io_in_5_Im(FFT_sr_v2_streaming_nrv_io_in_5_Im),
    .io_in_6_Re(FFT_sr_v2_streaming_nrv_io_in_6_Re),
    .io_in_6_Im(FFT_sr_v2_streaming_nrv_io_in_6_Im),
    .io_in_7_Re(FFT_sr_v2_streaming_nrv_io_in_7_Re),
    .io_in_7_Im(FFT_sr_v2_streaming_nrv_io_in_7_Im),
    .io_in_8_Re(FFT_sr_v2_streaming_nrv_io_in_8_Re),
    .io_in_8_Im(FFT_sr_v2_streaming_nrv_io_in_8_Im),
    .io_in_9_Re(FFT_sr_v2_streaming_nrv_io_in_9_Re),
    .io_in_9_Im(FFT_sr_v2_streaming_nrv_io_in_9_Im),
    .io_in_10_Re(FFT_sr_v2_streaming_nrv_io_in_10_Re),
    .io_in_10_Im(FFT_sr_v2_streaming_nrv_io_in_10_Im),
    .io_in_11_Re(FFT_sr_v2_streaming_nrv_io_in_11_Re),
    .io_in_11_Im(FFT_sr_v2_streaming_nrv_io_in_11_Im),
    .io_in_12_Re(FFT_sr_v2_streaming_nrv_io_in_12_Re),
    .io_in_12_Im(FFT_sr_v2_streaming_nrv_io_in_12_Im),
    .io_in_13_Re(FFT_sr_v2_streaming_nrv_io_in_13_Re),
    .io_in_13_Im(FFT_sr_v2_streaming_nrv_io_in_13_Im),
    .io_in_14_Re(FFT_sr_v2_streaming_nrv_io_in_14_Re),
    .io_in_14_Im(FFT_sr_v2_streaming_nrv_io_in_14_Im),
    .io_in_15_Re(FFT_sr_v2_streaming_nrv_io_in_15_Re),
    .io_in_15_Im(FFT_sr_v2_streaming_nrv_io_in_15_Im),
    .io_in_ready(FFT_sr_v2_streaming_nrv_io_in_ready),
    .io_out_0_Re(FFT_sr_v2_streaming_nrv_io_out_0_Re),
    .io_out_0_Im(FFT_sr_v2_streaming_nrv_io_out_0_Im),
    .io_out_1_Re(FFT_sr_v2_streaming_nrv_io_out_1_Re),
    .io_out_1_Im(FFT_sr_v2_streaming_nrv_io_out_1_Im),
    .io_out_2_Re(FFT_sr_v2_streaming_nrv_io_out_2_Re),
    .io_out_2_Im(FFT_sr_v2_streaming_nrv_io_out_2_Im),
    .io_out_3_Re(FFT_sr_v2_streaming_nrv_io_out_3_Re),
    .io_out_3_Im(FFT_sr_v2_streaming_nrv_io_out_3_Im),
    .io_out_4_Re(FFT_sr_v2_streaming_nrv_io_out_4_Re),
    .io_out_4_Im(FFT_sr_v2_streaming_nrv_io_out_4_Im),
    .io_out_5_Re(FFT_sr_v2_streaming_nrv_io_out_5_Re),
    .io_out_5_Im(FFT_sr_v2_streaming_nrv_io_out_5_Im),
    .io_out_6_Re(FFT_sr_v2_streaming_nrv_io_out_6_Re),
    .io_out_6_Im(FFT_sr_v2_streaming_nrv_io_out_6_Im),
    .io_out_7_Re(FFT_sr_v2_streaming_nrv_io_out_7_Re),
    .io_out_7_Im(FFT_sr_v2_streaming_nrv_io_out_7_Im),
    .io_out_8_Re(FFT_sr_v2_streaming_nrv_io_out_8_Re),
    .io_out_8_Im(FFT_sr_v2_streaming_nrv_io_out_8_Im),
    .io_out_9_Re(FFT_sr_v2_streaming_nrv_io_out_9_Re),
    .io_out_9_Im(FFT_sr_v2_streaming_nrv_io_out_9_Im),
    .io_out_10_Re(FFT_sr_v2_streaming_nrv_io_out_10_Re),
    .io_out_10_Im(FFT_sr_v2_streaming_nrv_io_out_10_Im),
    .io_out_11_Re(FFT_sr_v2_streaming_nrv_io_out_11_Re),
    .io_out_11_Im(FFT_sr_v2_streaming_nrv_io_out_11_Im),
    .io_out_12_Re(FFT_sr_v2_streaming_nrv_io_out_12_Re),
    .io_out_12_Im(FFT_sr_v2_streaming_nrv_io_out_12_Im),
    .io_out_13_Re(FFT_sr_v2_streaming_nrv_io_out_13_Re),
    .io_out_13_Im(FFT_sr_v2_streaming_nrv_io_out_13_Im),
    .io_out_14_Re(FFT_sr_v2_streaming_nrv_io_out_14_Re),
    .io_out_14_Im(FFT_sr_v2_streaming_nrv_io_out_14_Im),
    .io_out_15_Re(FFT_sr_v2_streaming_nrv_io_out_15_Re),
    .io_out_15_Im(FFT_sr_v2_streaming_nrv_io_out_15_Im)
  );
  DFT_r_v2_40 DFT_r_v2 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_clock),
    .reset(DFT_r_v2_reset),
    .io_in_0_Re(DFT_r_v2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_io_out_2_Im)
  );
  DFT_r_v2_40 DFT_r_v2_1 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_1_clock),
    .reset(DFT_r_v2_1_reset),
    .io_in_0_Re(DFT_r_v2_1_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_1_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_1_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_1_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_1_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_1_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_1_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_1_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_1_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_1_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_1_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_1_io_out_2_Im)
  );
  DFT_r_v2_40 DFT_r_v2_2 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_2_clock),
    .reset(DFT_r_v2_2_reset),
    .io_in_0_Re(DFT_r_v2_2_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_2_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_2_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_2_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_2_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_2_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_2_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_2_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_2_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_2_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_2_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_2_io_out_2_Im)
  );
  DFT_r_v2_40 DFT_r_v2_3 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_3_clock),
    .reset(DFT_r_v2_3_reset),
    .io_in_0_Re(DFT_r_v2_3_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_3_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_3_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_3_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_3_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_3_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_3_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_3_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_3_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_3_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_3_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_3_io_out_2_Im)
  );
  DFT_r_v2_40 DFT_r_v2_4 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_4_clock),
    .reset(DFT_r_v2_4_reset),
    .io_in_0_Re(DFT_r_v2_4_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_4_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_4_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_4_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_4_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_4_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_4_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_4_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_4_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_4_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_4_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_4_io_out_2_Im)
  );
  DFT_r_v2_40 DFT_r_v2_5 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_5_clock),
    .reset(DFT_r_v2_5_reset),
    .io_in_0_Re(DFT_r_v2_5_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_5_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_5_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_5_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_5_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_5_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_5_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_5_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_5_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_5_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_5_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_5_io_out_2_Im)
  );
  DFT_r_v2_40 DFT_r_v2_6 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_6_clock),
    .reset(DFT_r_v2_6_reset),
    .io_in_0_Re(DFT_r_v2_6_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_6_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_6_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_6_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_6_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_6_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_6_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_6_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_6_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_6_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_6_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_6_io_out_2_Im)
  );
  DFT_r_v2_40 DFT_r_v2_7 ( // @[FFTDesigns.scala 6457:32]
    .clock(DFT_r_v2_7_clock),
    .reset(DFT_r_v2_7_reset),
    .io_in_0_Re(DFT_r_v2_7_io_in_0_Re),
    .io_in_0_Im(DFT_r_v2_7_io_in_0_Im),
    .io_in_1_Re(DFT_r_v2_7_io_in_1_Re),
    .io_in_1_Im(DFT_r_v2_7_io_in_1_Im),
    .io_in_2_Re(DFT_r_v2_7_io_in_2_Re),
    .io_in_2_Im(DFT_r_v2_7_io_in_2_Im),
    .io_out_0_Re(DFT_r_v2_7_io_out_0_Re),
    .io_out_0_Im(DFT_r_v2_7_io_out_0_Im),
    .io_out_1_Re(DFT_r_v2_7_io_out_1_Re),
    .io_out_1_Im(DFT_r_v2_7_io_out_1_Im),
    .io_out_2_Re(DFT_r_v2_7_io_out_2_Re),
    .io_out_2_Im(DFT_r_v2_7_io_out_2_Im)
  );
  PermutationsWithStreaming_6 PermutationsWithStreaming ( // @[FFTDesigns.scala 6468:32]
    .clock(PermutationsWithStreaming_clock),
    .reset(PermutationsWithStreaming_reset),
    .io_in_0_Re(PermutationsWithStreaming_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_io_in_15_Im),
    .io_in_en_0(PermutationsWithStreaming_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_io_in_en_8),
    .io_in_en_9(PermutationsWithStreaming_io_in_en_9),
    .io_in_en_10(PermutationsWithStreaming_io_in_en_10),
    .io_in_en_11(PermutationsWithStreaming_io_in_en_11),
    .io_in_en_12(PermutationsWithStreaming_io_in_en_12),
    .io_out_0_Re(PermutationsWithStreaming_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_io_out_15_Im)
  );
  PermutationsWithStreaming_mr PermutationsWithStreaming_mr ( // @[FFTDesigns.scala 6469:32]
    .clock(PermutationsWithStreaming_mr_clock),
    .reset(PermutationsWithStreaming_mr_reset),
    .io_in_0_Re(PermutationsWithStreaming_mr_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_mr_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_mr_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_mr_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_mr_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_mr_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_mr_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_mr_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_mr_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_mr_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_mr_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_mr_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_mr_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_mr_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_mr_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_mr_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_mr_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_mr_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_mr_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_mr_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_mr_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_mr_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_mr_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_mr_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_mr_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_mr_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_mr_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_mr_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_mr_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_mr_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_mr_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_mr_io_in_15_Im),
    .io_in_en_0(PermutationsWithStreaming_mr_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_mr_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_mr_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_mr_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_mr_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_mr_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_mr_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_mr_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_mr_io_in_en_8),
    .io_in_en_9(PermutationsWithStreaming_mr_io_in_en_9),
    .io_in_en_10(PermutationsWithStreaming_mr_io_in_en_10),
    .io_in_en_11(PermutationsWithStreaming_mr_io_in_en_11),
    .io_in_en_12(PermutationsWithStreaming_mr_io_in_en_12),
    .io_out_0_Re(PermutationsWithStreaming_mr_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_mr_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_mr_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_mr_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_mr_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_mr_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_mr_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_mr_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_mr_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_mr_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_mr_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_mr_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_mr_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_mr_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_mr_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_mr_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_mr_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_mr_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_mr_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_mr_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_mr_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_mr_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_mr_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_mr_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_mr_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_mr_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_mr_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_mr_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_mr_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_mr_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_mr_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_mr_io_out_15_Im),
    .io_out_16_Re(PermutationsWithStreaming_mr_io_out_16_Re),
    .io_out_16_Im(PermutationsWithStreaming_mr_io_out_16_Im),
    .io_out_17_Re(PermutationsWithStreaming_mr_io_out_17_Re),
    .io_out_17_Im(PermutationsWithStreaming_mr_io_out_17_Im),
    .io_out_18_Re(PermutationsWithStreaming_mr_io_out_18_Re),
    .io_out_18_Im(PermutationsWithStreaming_mr_io_out_18_Im),
    .io_out_19_Re(PermutationsWithStreaming_mr_io_out_19_Re),
    .io_out_19_Im(PermutationsWithStreaming_mr_io_out_19_Im),
    .io_out_20_Re(PermutationsWithStreaming_mr_io_out_20_Re),
    .io_out_20_Im(PermutationsWithStreaming_mr_io_out_20_Im),
    .io_out_21_Re(PermutationsWithStreaming_mr_io_out_21_Re),
    .io_out_21_Im(PermutationsWithStreaming_mr_io_out_21_Im),
    .io_out_22_Re(PermutationsWithStreaming_mr_io_out_22_Re),
    .io_out_22_Im(PermutationsWithStreaming_mr_io_out_22_Im),
    .io_out_23_Re(PermutationsWithStreaming_mr_io_out_23_Re),
    .io_out_23_Im(PermutationsWithStreaming_mr_io_out_23_Im)
  );
  PermutationsWithStreaming_mr_1 PermutationsWithStreaming_mr_1 ( // @[FFTDesigns.scala 6470:32]
    .clock(PermutationsWithStreaming_mr_1_clock),
    .reset(PermutationsWithStreaming_mr_1_reset),
    .io_in_0_Re(PermutationsWithStreaming_mr_1_io_in_0_Re),
    .io_in_0_Im(PermutationsWithStreaming_mr_1_io_in_0_Im),
    .io_in_1_Re(PermutationsWithStreaming_mr_1_io_in_1_Re),
    .io_in_1_Im(PermutationsWithStreaming_mr_1_io_in_1_Im),
    .io_in_2_Re(PermutationsWithStreaming_mr_1_io_in_2_Re),
    .io_in_2_Im(PermutationsWithStreaming_mr_1_io_in_2_Im),
    .io_in_3_Re(PermutationsWithStreaming_mr_1_io_in_3_Re),
    .io_in_3_Im(PermutationsWithStreaming_mr_1_io_in_3_Im),
    .io_in_4_Re(PermutationsWithStreaming_mr_1_io_in_4_Re),
    .io_in_4_Im(PermutationsWithStreaming_mr_1_io_in_4_Im),
    .io_in_5_Re(PermutationsWithStreaming_mr_1_io_in_5_Re),
    .io_in_5_Im(PermutationsWithStreaming_mr_1_io_in_5_Im),
    .io_in_6_Re(PermutationsWithStreaming_mr_1_io_in_6_Re),
    .io_in_6_Im(PermutationsWithStreaming_mr_1_io_in_6_Im),
    .io_in_7_Re(PermutationsWithStreaming_mr_1_io_in_7_Re),
    .io_in_7_Im(PermutationsWithStreaming_mr_1_io_in_7_Im),
    .io_in_8_Re(PermutationsWithStreaming_mr_1_io_in_8_Re),
    .io_in_8_Im(PermutationsWithStreaming_mr_1_io_in_8_Im),
    .io_in_9_Re(PermutationsWithStreaming_mr_1_io_in_9_Re),
    .io_in_9_Im(PermutationsWithStreaming_mr_1_io_in_9_Im),
    .io_in_10_Re(PermutationsWithStreaming_mr_1_io_in_10_Re),
    .io_in_10_Im(PermutationsWithStreaming_mr_1_io_in_10_Im),
    .io_in_11_Re(PermutationsWithStreaming_mr_1_io_in_11_Re),
    .io_in_11_Im(PermutationsWithStreaming_mr_1_io_in_11_Im),
    .io_in_12_Re(PermutationsWithStreaming_mr_1_io_in_12_Re),
    .io_in_12_Im(PermutationsWithStreaming_mr_1_io_in_12_Im),
    .io_in_13_Re(PermutationsWithStreaming_mr_1_io_in_13_Re),
    .io_in_13_Im(PermutationsWithStreaming_mr_1_io_in_13_Im),
    .io_in_14_Re(PermutationsWithStreaming_mr_1_io_in_14_Re),
    .io_in_14_Im(PermutationsWithStreaming_mr_1_io_in_14_Im),
    .io_in_15_Re(PermutationsWithStreaming_mr_1_io_in_15_Re),
    .io_in_15_Im(PermutationsWithStreaming_mr_1_io_in_15_Im),
    .io_in_16_Re(PermutationsWithStreaming_mr_1_io_in_16_Re),
    .io_in_16_Im(PermutationsWithStreaming_mr_1_io_in_16_Im),
    .io_in_17_Re(PermutationsWithStreaming_mr_1_io_in_17_Re),
    .io_in_17_Im(PermutationsWithStreaming_mr_1_io_in_17_Im),
    .io_in_18_Re(PermutationsWithStreaming_mr_1_io_in_18_Re),
    .io_in_18_Im(PermutationsWithStreaming_mr_1_io_in_18_Im),
    .io_in_19_Re(PermutationsWithStreaming_mr_1_io_in_19_Re),
    .io_in_19_Im(PermutationsWithStreaming_mr_1_io_in_19_Im),
    .io_in_20_Re(PermutationsWithStreaming_mr_1_io_in_20_Re),
    .io_in_20_Im(PermutationsWithStreaming_mr_1_io_in_20_Im),
    .io_in_21_Re(PermutationsWithStreaming_mr_1_io_in_21_Re),
    .io_in_21_Im(PermutationsWithStreaming_mr_1_io_in_21_Im),
    .io_in_22_Re(PermutationsWithStreaming_mr_1_io_in_22_Re),
    .io_in_22_Im(PermutationsWithStreaming_mr_1_io_in_22_Im),
    .io_in_23_Re(PermutationsWithStreaming_mr_1_io_in_23_Re),
    .io_in_23_Im(PermutationsWithStreaming_mr_1_io_in_23_Im),
    .io_in_en_0(PermutationsWithStreaming_mr_1_io_in_en_0),
    .io_in_en_1(PermutationsWithStreaming_mr_1_io_in_en_1),
    .io_in_en_2(PermutationsWithStreaming_mr_1_io_in_en_2),
    .io_in_en_3(PermutationsWithStreaming_mr_1_io_in_en_3),
    .io_in_en_4(PermutationsWithStreaming_mr_1_io_in_en_4),
    .io_in_en_5(PermutationsWithStreaming_mr_1_io_in_en_5),
    .io_in_en_6(PermutationsWithStreaming_mr_1_io_in_en_6),
    .io_in_en_7(PermutationsWithStreaming_mr_1_io_in_en_7),
    .io_in_en_8(PermutationsWithStreaming_mr_1_io_in_en_8),
    .io_in_en_9(PermutationsWithStreaming_mr_1_io_in_en_9),
    .io_in_en_10(PermutationsWithStreaming_mr_1_io_in_en_10),
    .io_in_en_11(PermutationsWithStreaming_mr_1_io_in_en_11),
    .io_in_en_12(PermutationsWithStreaming_mr_1_io_in_en_12),
    .io_out_0_Re(PermutationsWithStreaming_mr_1_io_out_0_Re),
    .io_out_0_Im(PermutationsWithStreaming_mr_1_io_out_0_Im),
    .io_out_1_Re(PermutationsWithStreaming_mr_1_io_out_1_Re),
    .io_out_1_Im(PermutationsWithStreaming_mr_1_io_out_1_Im),
    .io_out_2_Re(PermutationsWithStreaming_mr_1_io_out_2_Re),
    .io_out_2_Im(PermutationsWithStreaming_mr_1_io_out_2_Im),
    .io_out_3_Re(PermutationsWithStreaming_mr_1_io_out_3_Re),
    .io_out_3_Im(PermutationsWithStreaming_mr_1_io_out_3_Im),
    .io_out_4_Re(PermutationsWithStreaming_mr_1_io_out_4_Re),
    .io_out_4_Im(PermutationsWithStreaming_mr_1_io_out_4_Im),
    .io_out_5_Re(PermutationsWithStreaming_mr_1_io_out_5_Re),
    .io_out_5_Im(PermutationsWithStreaming_mr_1_io_out_5_Im),
    .io_out_6_Re(PermutationsWithStreaming_mr_1_io_out_6_Re),
    .io_out_6_Im(PermutationsWithStreaming_mr_1_io_out_6_Im),
    .io_out_7_Re(PermutationsWithStreaming_mr_1_io_out_7_Re),
    .io_out_7_Im(PermutationsWithStreaming_mr_1_io_out_7_Im),
    .io_out_8_Re(PermutationsWithStreaming_mr_1_io_out_8_Re),
    .io_out_8_Im(PermutationsWithStreaming_mr_1_io_out_8_Im),
    .io_out_9_Re(PermutationsWithStreaming_mr_1_io_out_9_Re),
    .io_out_9_Im(PermutationsWithStreaming_mr_1_io_out_9_Im),
    .io_out_10_Re(PermutationsWithStreaming_mr_1_io_out_10_Re),
    .io_out_10_Im(PermutationsWithStreaming_mr_1_io_out_10_Im),
    .io_out_11_Re(PermutationsWithStreaming_mr_1_io_out_11_Re),
    .io_out_11_Im(PermutationsWithStreaming_mr_1_io_out_11_Im),
    .io_out_12_Re(PermutationsWithStreaming_mr_1_io_out_12_Re),
    .io_out_12_Im(PermutationsWithStreaming_mr_1_io_out_12_Im),
    .io_out_13_Re(PermutationsWithStreaming_mr_1_io_out_13_Re),
    .io_out_13_Im(PermutationsWithStreaming_mr_1_io_out_13_Im),
    .io_out_14_Re(PermutationsWithStreaming_mr_1_io_out_14_Re),
    .io_out_14_Im(PermutationsWithStreaming_mr_1_io_out_14_Im),
    .io_out_15_Re(PermutationsWithStreaming_mr_1_io_out_15_Re),
    .io_out_15_Im(PermutationsWithStreaming_mr_1_io_out_15_Im)
  );
  TwiddleFactorsStreamed_mr_v2 TwiddleFactorsStreamed_mr_v2 ( // @[FFTDesigns.scala 6471:32]
    .clock(TwiddleFactorsStreamed_mr_v2_clock),
    .reset(TwiddleFactorsStreamed_mr_v2_reset),
    .io_in_0_Re(TwiddleFactorsStreamed_mr_v2_io_in_0_Re),
    .io_in_0_Im(TwiddleFactorsStreamed_mr_v2_io_in_0_Im),
    .io_in_1_Re(TwiddleFactorsStreamed_mr_v2_io_in_1_Re),
    .io_in_1_Im(TwiddleFactorsStreamed_mr_v2_io_in_1_Im),
    .io_in_2_Re(TwiddleFactorsStreamed_mr_v2_io_in_2_Re),
    .io_in_2_Im(TwiddleFactorsStreamed_mr_v2_io_in_2_Im),
    .io_in_3_Re(TwiddleFactorsStreamed_mr_v2_io_in_3_Re),
    .io_in_3_Im(TwiddleFactorsStreamed_mr_v2_io_in_3_Im),
    .io_in_4_Re(TwiddleFactorsStreamed_mr_v2_io_in_4_Re),
    .io_in_4_Im(TwiddleFactorsStreamed_mr_v2_io_in_4_Im),
    .io_in_5_Re(TwiddleFactorsStreamed_mr_v2_io_in_5_Re),
    .io_in_5_Im(TwiddleFactorsStreamed_mr_v2_io_in_5_Im),
    .io_in_6_Re(TwiddleFactorsStreamed_mr_v2_io_in_6_Re),
    .io_in_6_Im(TwiddleFactorsStreamed_mr_v2_io_in_6_Im),
    .io_in_7_Re(TwiddleFactorsStreamed_mr_v2_io_in_7_Re),
    .io_in_7_Im(TwiddleFactorsStreamed_mr_v2_io_in_7_Im),
    .io_in_8_Re(TwiddleFactorsStreamed_mr_v2_io_in_8_Re),
    .io_in_8_Im(TwiddleFactorsStreamed_mr_v2_io_in_8_Im),
    .io_in_9_Re(TwiddleFactorsStreamed_mr_v2_io_in_9_Re),
    .io_in_9_Im(TwiddleFactorsStreamed_mr_v2_io_in_9_Im),
    .io_in_10_Re(TwiddleFactorsStreamed_mr_v2_io_in_10_Re),
    .io_in_10_Im(TwiddleFactorsStreamed_mr_v2_io_in_10_Im),
    .io_in_11_Re(TwiddleFactorsStreamed_mr_v2_io_in_11_Re),
    .io_in_11_Im(TwiddleFactorsStreamed_mr_v2_io_in_11_Im),
    .io_in_12_Re(TwiddleFactorsStreamed_mr_v2_io_in_12_Re),
    .io_in_12_Im(TwiddleFactorsStreamed_mr_v2_io_in_12_Im),
    .io_in_13_Re(TwiddleFactorsStreamed_mr_v2_io_in_13_Re),
    .io_in_13_Im(TwiddleFactorsStreamed_mr_v2_io_in_13_Im),
    .io_in_14_Re(TwiddleFactorsStreamed_mr_v2_io_in_14_Re),
    .io_in_14_Im(TwiddleFactorsStreamed_mr_v2_io_in_14_Im),
    .io_in_15_Re(TwiddleFactorsStreamed_mr_v2_io_in_15_Re),
    .io_in_15_Im(TwiddleFactorsStreamed_mr_v2_io_in_15_Im),
    .io_in_16_Re(TwiddleFactorsStreamed_mr_v2_io_in_16_Re),
    .io_in_16_Im(TwiddleFactorsStreamed_mr_v2_io_in_16_Im),
    .io_in_17_Re(TwiddleFactorsStreamed_mr_v2_io_in_17_Re),
    .io_in_17_Im(TwiddleFactorsStreamed_mr_v2_io_in_17_Im),
    .io_in_18_Re(TwiddleFactorsStreamed_mr_v2_io_in_18_Re),
    .io_in_18_Im(TwiddleFactorsStreamed_mr_v2_io_in_18_Im),
    .io_in_19_Re(TwiddleFactorsStreamed_mr_v2_io_in_19_Re),
    .io_in_19_Im(TwiddleFactorsStreamed_mr_v2_io_in_19_Im),
    .io_in_20_Re(TwiddleFactorsStreamed_mr_v2_io_in_20_Re),
    .io_in_20_Im(TwiddleFactorsStreamed_mr_v2_io_in_20_Im),
    .io_in_21_Re(TwiddleFactorsStreamed_mr_v2_io_in_21_Re),
    .io_in_21_Im(TwiddleFactorsStreamed_mr_v2_io_in_21_Im),
    .io_in_22_Re(TwiddleFactorsStreamed_mr_v2_io_in_22_Re),
    .io_in_22_Im(TwiddleFactorsStreamed_mr_v2_io_in_22_Im),
    .io_in_23_Re(TwiddleFactorsStreamed_mr_v2_io_in_23_Re),
    .io_in_23_Im(TwiddleFactorsStreamed_mr_v2_io_in_23_Im),
    .io_in_en_0(TwiddleFactorsStreamed_mr_v2_io_in_en_0),
    .io_in_en_1(TwiddleFactorsStreamed_mr_v2_io_in_en_1),
    .io_out_0_Re(TwiddleFactorsStreamed_mr_v2_io_out_0_Re),
    .io_out_0_Im(TwiddleFactorsStreamed_mr_v2_io_out_0_Im),
    .io_out_1_Re(TwiddleFactorsStreamed_mr_v2_io_out_1_Re),
    .io_out_1_Im(TwiddleFactorsStreamed_mr_v2_io_out_1_Im),
    .io_out_2_Re(TwiddleFactorsStreamed_mr_v2_io_out_2_Re),
    .io_out_2_Im(TwiddleFactorsStreamed_mr_v2_io_out_2_Im),
    .io_out_3_Re(TwiddleFactorsStreamed_mr_v2_io_out_3_Re),
    .io_out_3_Im(TwiddleFactorsStreamed_mr_v2_io_out_3_Im),
    .io_out_4_Re(TwiddleFactorsStreamed_mr_v2_io_out_4_Re),
    .io_out_4_Im(TwiddleFactorsStreamed_mr_v2_io_out_4_Im),
    .io_out_5_Re(TwiddleFactorsStreamed_mr_v2_io_out_5_Re),
    .io_out_5_Im(TwiddleFactorsStreamed_mr_v2_io_out_5_Im),
    .io_out_6_Re(TwiddleFactorsStreamed_mr_v2_io_out_6_Re),
    .io_out_6_Im(TwiddleFactorsStreamed_mr_v2_io_out_6_Im),
    .io_out_7_Re(TwiddleFactorsStreamed_mr_v2_io_out_7_Re),
    .io_out_7_Im(TwiddleFactorsStreamed_mr_v2_io_out_7_Im),
    .io_out_8_Re(TwiddleFactorsStreamed_mr_v2_io_out_8_Re),
    .io_out_8_Im(TwiddleFactorsStreamed_mr_v2_io_out_8_Im),
    .io_out_9_Re(TwiddleFactorsStreamed_mr_v2_io_out_9_Re),
    .io_out_9_Im(TwiddleFactorsStreamed_mr_v2_io_out_9_Im),
    .io_out_10_Re(TwiddleFactorsStreamed_mr_v2_io_out_10_Re),
    .io_out_10_Im(TwiddleFactorsStreamed_mr_v2_io_out_10_Im),
    .io_out_11_Re(TwiddleFactorsStreamed_mr_v2_io_out_11_Re),
    .io_out_11_Im(TwiddleFactorsStreamed_mr_v2_io_out_11_Im),
    .io_out_12_Re(TwiddleFactorsStreamed_mr_v2_io_out_12_Re),
    .io_out_12_Im(TwiddleFactorsStreamed_mr_v2_io_out_12_Im),
    .io_out_13_Re(TwiddleFactorsStreamed_mr_v2_io_out_13_Re),
    .io_out_13_Im(TwiddleFactorsStreamed_mr_v2_io_out_13_Im),
    .io_out_14_Re(TwiddleFactorsStreamed_mr_v2_io_out_14_Re),
    .io_out_14_Im(TwiddleFactorsStreamed_mr_v2_io_out_14_Im),
    .io_out_15_Re(TwiddleFactorsStreamed_mr_v2_io_out_15_Re),
    .io_out_15_Im(TwiddleFactorsStreamed_mr_v2_io_out_15_Im),
    .io_out_16_Re(TwiddleFactorsStreamed_mr_v2_io_out_16_Re),
    .io_out_16_Im(TwiddleFactorsStreamed_mr_v2_io_out_16_Im),
    .io_out_17_Re(TwiddleFactorsStreamed_mr_v2_io_out_17_Re),
    .io_out_17_Im(TwiddleFactorsStreamed_mr_v2_io_out_17_Im),
    .io_out_18_Re(TwiddleFactorsStreamed_mr_v2_io_out_18_Re),
    .io_out_18_Im(TwiddleFactorsStreamed_mr_v2_io_out_18_Im),
    .io_out_19_Re(TwiddleFactorsStreamed_mr_v2_io_out_19_Re),
    .io_out_19_Im(TwiddleFactorsStreamed_mr_v2_io_out_19_Im),
    .io_out_20_Re(TwiddleFactorsStreamed_mr_v2_io_out_20_Re),
    .io_out_20_Im(TwiddleFactorsStreamed_mr_v2_io_out_20_Im),
    .io_out_21_Re(TwiddleFactorsStreamed_mr_v2_io_out_21_Re),
    .io_out_21_Im(TwiddleFactorsStreamed_mr_v2_io_out_21_Im),
    .io_out_22_Re(TwiddleFactorsStreamed_mr_v2_io_out_22_Re),
    .io_out_22_Im(TwiddleFactorsStreamed_mr_v2_io_out_22_Im),
    .io_out_23_Re(TwiddleFactorsStreamed_mr_v2_io_out_23_Re),
    .io_out_23_Im(TwiddleFactorsStreamed_mr_v2_io_out_23_Im)
  );
  assign io_out_validate = out_regdelay; // @[FFTDesigns.scala 6560:23]
  assign io_out_0_Re = results_0_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_0_Im = results_0_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_1_Re = results_1_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_1_Im = results_1_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_2_Re = results_2_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_2_Im = results_2_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_3_Re = results_3_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_3_Im = results_3_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_4_Re = results_4_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_4_Im = results_4_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_5_Re = results_5_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_5_Im = results_5_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_6_Re = results_6_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_6_Im = results_6_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_7_Re = results_7_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_7_Im = results_7_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_8_Re = results_8_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_8_Im = results_8_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_9_Re = results_9_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_9_Im = results_9_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_10_Re = results_10_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_10_Im = results_10_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_11_Re = results_11_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_11_Im = results_11_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_12_Re = results_12_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_12_Im = results_12_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_13_Re = results_13_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_13_Im = results_13_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_14_Re = results_14_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_14_Im = results_14_Im; // @[FFTDesigns.scala 6561:14]
  assign io_out_15_Re = results_15_Re; // @[FFTDesigns.scala 6561:14]
  assign io_out_15_Im = results_15_Im; // @[FFTDesigns.scala 6561:14]
  assign FFT_sr_v2_streaming_nrv_clock = clock;
  assign FFT_sr_v2_streaming_nrv_reset = reset;
  assign FFT_sr_v2_streaming_nrv_io_in_0_Re = PermutationsWithStreaming_io_out_0_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_0_Im = PermutationsWithStreaming_io_out_0_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_1_Re = PermutationsWithStreaming_io_out_1_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_1_Im = PermutationsWithStreaming_io_out_1_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_2_Re = PermutationsWithStreaming_io_out_2_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_2_Im = PermutationsWithStreaming_io_out_2_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_3_Re = PermutationsWithStreaming_io_out_3_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_3_Im = PermutationsWithStreaming_io_out_3_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_4_Re = PermutationsWithStreaming_io_out_4_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_4_Im = PermutationsWithStreaming_io_out_4_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_5_Re = PermutationsWithStreaming_io_out_5_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_5_Im = PermutationsWithStreaming_io_out_5_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_6_Re = PermutationsWithStreaming_io_out_6_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_6_Im = PermutationsWithStreaming_io_out_6_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_7_Re = PermutationsWithStreaming_io_out_7_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_7_Im = PermutationsWithStreaming_io_out_7_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_8_Re = PermutationsWithStreaming_io_out_8_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_8_Im = PermutationsWithStreaming_io_out_8_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_9_Re = PermutationsWithStreaming_io_out_9_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_9_Im = PermutationsWithStreaming_io_out_9_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_10_Re = PermutationsWithStreaming_io_out_10_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_10_Im = PermutationsWithStreaming_io_out_10_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_11_Re = PermutationsWithStreaming_io_out_11_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_11_Im = PermutationsWithStreaming_io_out_11_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_12_Re = PermutationsWithStreaming_io_out_12_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_12_Im = PermutationsWithStreaming_io_out_12_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_13_Re = PermutationsWithStreaming_io_out_13_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_13_Im = PermutationsWithStreaming_io_out_13_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_14_Re = PermutationsWithStreaming_io_out_14_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_14_Im = PermutationsWithStreaming_io_out_14_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_15_Re = PermutationsWithStreaming_io_out_15_Re; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_15_Im = PermutationsWithStreaming_io_out_15_Im; // @[FFTDesigns.scala 6535:27]
  assign FFT_sr_v2_streaming_nrv_io_in_ready = Perm_regdelays1_0_11; // @[FFTDesigns.scala 6536:33]
  assign DFT_r_v2_clock = clock;
  assign DFT_r_v2_reset = reset;
  assign DFT_r_v2_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_0_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_0_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_1_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_1_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_2_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_2_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_clock = clock;
  assign DFT_r_v2_1_reset = reset;
  assign DFT_r_v2_1_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_3_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_3_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_4_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_4_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_5_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_1_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_5_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_clock = clock;
  assign DFT_r_v2_2_reset = reset;
  assign DFT_r_v2_2_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_6_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_6_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_7_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_7_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_8_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_2_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_8_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_clock = clock;
  assign DFT_r_v2_3_reset = reset;
  assign DFT_r_v2_3_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_9_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_9_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_10_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_10_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_11_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_3_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_11_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_4_clock = clock;
  assign DFT_r_v2_4_reset = reset;
  assign DFT_r_v2_4_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_12_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_4_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_12_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_4_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_13_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_4_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_13_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_4_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_14_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_4_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_14_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_5_clock = clock;
  assign DFT_r_v2_5_reset = reset;
  assign DFT_r_v2_5_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_15_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_5_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_15_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_5_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_16_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_5_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_16_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_5_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_17_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_5_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_17_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_6_clock = clock;
  assign DFT_r_v2_6_reset = reset;
  assign DFT_r_v2_6_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_18_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_6_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_18_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_6_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_19_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_6_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_19_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_6_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_20_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_6_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_20_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_7_clock = clock;
  assign DFT_r_v2_7_reset = reset;
  assign DFT_r_v2_7_io_in_0_Re = TwiddleFactorsStreamed_mr_v2_io_out_21_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_7_io_in_0_Im = TwiddleFactorsStreamed_mr_v2_io_out_21_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_7_io_in_1_Re = TwiddleFactorsStreamed_mr_v2_io_out_22_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_7_io_in_1_Im = TwiddleFactorsStreamed_mr_v2_io_out_22_Im; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_7_io_in_2_Re = TwiddleFactorsStreamed_mr_v2_io_out_23_Re; // @[FFTDesigns.scala 6547:37]
  assign DFT_r_v2_7_io_in_2_Im = TwiddleFactorsStreamed_mr_v2_io_out_23_Im; // @[FFTDesigns.scala 6547:37]
  assign PermutationsWithStreaming_clock = clock;
  assign PermutationsWithStreaming_reset = reset;
  assign PermutationsWithStreaming_io_in_0_Re = io_in_0_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_0_Im = io_in_0_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_1_Re = io_in_1_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_1_Im = io_in_1_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_2_Re = io_in_2_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_2_Im = io_in_2_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_3_Re = io_in_3_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_3_Im = io_in_3_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_4_Re = io_in_4_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_4_Im = io_in_4_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_5_Re = io_in_5_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_5_Im = io_in_5_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_6_Re = io_in_6_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_6_Im = io_in_6_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_7_Re = io_in_7_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_7_Im = io_in_7_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_8_Re = io_in_8_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_8_Im = io_in_8_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_9_Re = io_in_9_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_9_Im = io_in_9_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_10_Re = io_in_10_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_10_Im = io_in_10_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_11_Re = io_in_11_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_11_Im = io_in_11_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_12_Re = io_in_12_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_12_Im = io_in_12_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_13_Re = io_in_13_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_13_Im = io_in_13_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_14_Re = io_in_14_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_14_Im = io_in_14_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_15_Re = io_in_15_Re; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_15_Im = io_in_15_Im; // @[FFTDesigns.scala 6486:31]
  assign PermutationsWithStreaming_io_in_en_0 = io_in_ready; // @[FFTDesigns.scala 6485:37]
  assign PermutationsWithStreaming_io_in_en_1 = Perm_regdelays1_0_0; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_2 = Perm_regdelays1_0_1; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_3 = Perm_regdelays1_0_2; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_4 = Perm_regdelays1_0_3; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_5 = Perm_regdelays1_0_4; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_6 = Perm_regdelays1_0_5; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_7 = Perm_regdelays1_0_6; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_8 = Perm_regdelays1_0_7; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_9 = Perm_regdelays1_0_8; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_10 = Perm_regdelays1_0_9; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_11 = Perm_regdelays1_0_10; // @[FFTDesigns.scala 6503:37]
  assign PermutationsWithStreaming_io_in_en_12 = Perm_regdelays1_0_11; // @[FFTDesigns.scala 6511:51]
  assign PermutationsWithStreaming_mr_clock = clock;
  assign PermutationsWithStreaming_mr_reset = reset;
  assign PermutationsWithStreaming_mr_io_in_0_Re = FFT_sr_v2_streaming_nrv_io_out_0_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_0_Im = FFT_sr_v2_streaming_nrv_io_out_0_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_1_Re = FFT_sr_v2_streaming_nrv_io_out_1_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_1_Im = FFT_sr_v2_streaming_nrv_io_out_1_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_2_Re = FFT_sr_v2_streaming_nrv_io_out_2_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_2_Im = FFT_sr_v2_streaming_nrv_io_out_2_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_3_Re = FFT_sr_v2_streaming_nrv_io_out_3_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_3_Im = FFT_sr_v2_streaming_nrv_io_out_3_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_4_Re = FFT_sr_v2_streaming_nrv_io_out_4_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_4_Im = FFT_sr_v2_streaming_nrv_io_out_4_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_5_Re = FFT_sr_v2_streaming_nrv_io_out_5_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_5_Im = FFT_sr_v2_streaming_nrv_io_out_5_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_6_Re = FFT_sr_v2_streaming_nrv_io_out_6_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_6_Im = FFT_sr_v2_streaming_nrv_io_out_6_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_7_Re = FFT_sr_v2_streaming_nrv_io_out_7_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_7_Im = FFT_sr_v2_streaming_nrv_io_out_7_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_8_Re = FFT_sr_v2_streaming_nrv_io_out_8_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_8_Im = FFT_sr_v2_streaming_nrv_io_out_8_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_9_Re = FFT_sr_v2_streaming_nrv_io_out_9_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_9_Im = FFT_sr_v2_streaming_nrv_io_out_9_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_10_Re = FFT_sr_v2_streaming_nrv_io_out_10_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_10_Im = FFT_sr_v2_streaming_nrv_io_out_10_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_11_Re = FFT_sr_v2_streaming_nrv_io_out_11_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_11_Im = FFT_sr_v2_streaming_nrv_io_out_11_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_12_Re = FFT_sr_v2_streaming_nrv_io_out_12_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_12_Im = FFT_sr_v2_streaming_nrv_io_out_12_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_13_Re = FFT_sr_v2_streaming_nrv_io_out_13_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_13_Im = FFT_sr_v2_streaming_nrv_io_out_13_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_14_Re = FFT_sr_v2_streaming_nrv_io_out_14_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_14_Im = FFT_sr_v2_streaming_nrv_io_out_14_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_15_Re = FFT_sr_v2_streaming_nrv_io_out_15_Re; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_15_Im = FFT_sr_v2_streaming_nrv_io_out_15_Im; // @[FFTDesigns.scala 6490:31]
  assign PermutationsWithStreaming_mr_io_in_en_0 = DFT_regdelays1_36; // @[FFTDesigns.scala 6489:37]
  assign PermutationsWithStreaming_mr_io_in_en_1 = Perm_regdelays1_1_0; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_2 = Perm_regdelays1_1_1; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_3 = Perm_regdelays1_1_2; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_4 = Perm_regdelays1_1_3; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_5 = Perm_regdelays1_1_4; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_6 = Perm_regdelays1_1_5; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_7 = Perm_regdelays1_1_6; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_8 = Perm_regdelays1_1_7; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_9 = Perm_regdelays1_1_8; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_10 = Perm_regdelays1_1_9; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_11 = Perm_regdelays1_1_10; // @[FFTDesigns.scala 6505:37]
  assign PermutationsWithStreaming_mr_io_in_en_12 = Perm_regdelays1_1_11; // @[FFTDesigns.scala 6513:51]
  assign PermutationsWithStreaming_mr_1_clock = clock;
  assign PermutationsWithStreaming_mr_1_reset = reset;
  assign PermutationsWithStreaming_mr_1_io_in_0_Re = DFT_r_v2_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_0_Im = DFT_r_v2_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_1_Re = DFT_r_v2_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_1_Im = DFT_r_v2_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_2_Re = DFT_r_v2_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_2_Im = DFT_r_v2_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_3_Re = DFT_r_v2_1_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_3_Im = DFT_r_v2_1_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_4_Re = DFT_r_v2_1_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_4_Im = DFT_r_v2_1_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_5_Re = DFT_r_v2_1_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_5_Im = DFT_r_v2_1_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_6_Re = DFT_r_v2_2_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_6_Im = DFT_r_v2_2_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_7_Re = DFT_r_v2_2_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_7_Im = DFT_r_v2_2_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_8_Re = DFT_r_v2_2_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_8_Im = DFT_r_v2_2_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_9_Re = DFT_r_v2_3_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_9_Im = DFT_r_v2_3_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_10_Re = DFT_r_v2_3_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_10_Im = DFT_r_v2_3_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_11_Re = DFT_r_v2_3_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_11_Im = DFT_r_v2_3_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_12_Re = DFT_r_v2_4_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_12_Im = DFT_r_v2_4_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_13_Re = DFT_r_v2_4_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_13_Im = DFT_r_v2_4_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_14_Re = DFT_r_v2_4_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_14_Im = DFT_r_v2_4_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_15_Re = DFT_r_v2_5_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_15_Im = DFT_r_v2_5_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_16_Re = DFT_r_v2_5_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_16_Im = DFT_r_v2_5_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_17_Re = DFT_r_v2_5_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_17_Im = DFT_r_v2_5_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_18_Re = DFT_r_v2_6_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_18_Im = DFT_r_v2_6_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_19_Re = DFT_r_v2_6_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_19_Im = DFT_r_v2_6_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_20_Re = DFT_r_v2_6_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_20_Im = DFT_r_v2_6_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_21_Re = DFT_r_v2_7_io_out_0_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_21_Im = DFT_r_v2_7_io_out_0_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_22_Re = DFT_r_v2_7_io_out_1_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_22_Im = DFT_r_v2_7_io_out_1_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_23_Re = DFT_r_v2_7_io_out_2_Re; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_23_Im = DFT_r_v2_7_io_out_2_Im; // @[FFTDesigns.scala 6496:45]
  assign PermutationsWithStreaming_mr_1_io_in_en_0 = DFT_regdelays2_3; // @[FFTDesigns.scala 6493:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_1 = Perm_regdelays1_2_0; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_2 = Perm_regdelays1_2_1; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_3 = Perm_regdelays1_2_2; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_4 = Perm_regdelays1_2_3; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_5 = Perm_regdelays1_2_4; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_6 = Perm_regdelays1_2_5; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_7 = Perm_regdelays1_2_6; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_8 = Perm_regdelays1_2_7; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_9 = Perm_regdelays1_2_8; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_10 = Perm_regdelays1_2_9; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_11 = Perm_regdelays1_2_10; // @[FFTDesigns.scala 6507:37]
  assign PermutationsWithStreaming_mr_1_io_in_en_12 = Perm_regdelays1_2_11; // @[FFTDesigns.scala 6515:51]
  assign TwiddleFactorsStreamed_mr_v2_clock = clock;
  assign TwiddleFactorsStreamed_mr_v2_reset = reset;
  assign TwiddleFactorsStreamed_mr_v2_io_in_0_Re = PermutationsWithStreaming_mr_io_out_0_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_0_Im = PermutationsWithStreaming_mr_io_out_0_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_1_Re = PermutationsWithStreaming_mr_io_out_1_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_1_Im = PermutationsWithStreaming_mr_io_out_1_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_2_Re = PermutationsWithStreaming_mr_io_out_2_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_2_Im = PermutationsWithStreaming_mr_io_out_2_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_3_Re = PermutationsWithStreaming_mr_io_out_3_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_3_Im = PermutationsWithStreaming_mr_io_out_3_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_4_Re = PermutationsWithStreaming_mr_io_out_4_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_4_Im = PermutationsWithStreaming_mr_io_out_4_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_5_Re = PermutationsWithStreaming_mr_io_out_5_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_5_Im = PermutationsWithStreaming_mr_io_out_5_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_6_Re = PermutationsWithStreaming_mr_io_out_6_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_6_Im = PermutationsWithStreaming_mr_io_out_6_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_7_Re = PermutationsWithStreaming_mr_io_out_7_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_7_Im = PermutationsWithStreaming_mr_io_out_7_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_8_Re = PermutationsWithStreaming_mr_io_out_8_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_8_Im = PermutationsWithStreaming_mr_io_out_8_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_9_Re = PermutationsWithStreaming_mr_io_out_9_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_9_Im = PermutationsWithStreaming_mr_io_out_9_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_10_Re = PermutationsWithStreaming_mr_io_out_10_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_10_Im = PermutationsWithStreaming_mr_io_out_10_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_11_Re = PermutationsWithStreaming_mr_io_out_11_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_11_Im = PermutationsWithStreaming_mr_io_out_11_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_12_Re = PermutationsWithStreaming_mr_io_out_12_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_12_Im = PermutationsWithStreaming_mr_io_out_12_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_13_Re = PermutationsWithStreaming_mr_io_out_13_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_13_Im = PermutationsWithStreaming_mr_io_out_13_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_14_Re = PermutationsWithStreaming_mr_io_out_14_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_14_Im = PermutationsWithStreaming_mr_io_out_14_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_15_Re = PermutationsWithStreaming_mr_io_out_15_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_15_Im = PermutationsWithStreaming_mr_io_out_15_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_16_Re = PermutationsWithStreaming_mr_io_out_16_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_16_Im = PermutationsWithStreaming_mr_io_out_16_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_17_Re = PermutationsWithStreaming_mr_io_out_17_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_17_Im = PermutationsWithStreaming_mr_io_out_17_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_18_Re = PermutationsWithStreaming_mr_io_out_18_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_18_Im = PermutationsWithStreaming_mr_io_out_18_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_19_Re = PermutationsWithStreaming_mr_io_out_19_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_19_Im = PermutationsWithStreaming_mr_io_out_19_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_20_Re = PermutationsWithStreaming_mr_io_out_20_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_20_Im = PermutationsWithStreaming_mr_io_out_20_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_21_Re = PermutationsWithStreaming_mr_io_out_21_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_21_Im = PermutationsWithStreaming_mr_io_out_21_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_22_Re = PermutationsWithStreaming_mr_io_out_22_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_22_Im = PermutationsWithStreaming_mr_io_out_22_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_23_Re = PermutationsWithStreaming_mr_io_out_23_Re; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_23_Im = PermutationsWithStreaming_mr_io_out_23_Im; // @[FFTDesigns.scala 6525:27]
  assign TwiddleFactorsStreamed_mr_v2_io_in_en_0 = Perm_regdelays1_1_11; // @[FFTDesigns.scala 6524:33]
  assign TwiddleFactorsStreamed_mr_v2_io_in_en_1 = Twid_regdelays_0; // @[FFTDesigns.scala 6528:33]
  always @(posedge clock) begin
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_0 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_0 <= Perm_regdelays1_0_11; // @[FFTDesigns.scala 6534:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_1 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_1 <= DFT_regdelays1_0; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_2 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_2 <= DFT_regdelays1_1; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_3 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_3 <= DFT_regdelays1_2; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_4 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_4 <= DFT_regdelays1_3; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_5 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_5 <= DFT_regdelays1_4; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_6 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_6 <= DFT_regdelays1_5; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_7 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_7 <= DFT_regdelays1_6; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_8 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_8 <= DFT_regdelays1_7; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_9 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_9 <= DFT_regdelays1_8; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_10 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_10 <= DFT_regdelays1_9; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_11 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_11 <= DFT_regdelays1_10; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_12 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_12 <= DFT_regdelays1_11; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_13 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_13 <= DFT_regdelays1_12; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_14 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_14 <= DFT_regdelays1_13; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_15 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_15 <= DFT_regdelays1_14; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_16 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_16 <= DFT_regdelays1_15; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_17 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_17 <= DFT_regdelays1_16; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_18 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_18 <= DFT_regdelays1_17; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_19 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_19 <= DFT_regdelays1_18; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_20 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_20 <= DFT_regdelays1_19; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_21 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_21 <= DFT_regdelays1_20; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_22 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_22 <= DFT_regdelays1_21; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_23 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_23 <= DFT_regdelays1_22; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_24 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_24 <= DFT_regdelays1_23; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_25 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_25 <= DFT_regdelays1_24; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_26 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_26 <= DFT_regdelays1_25; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_27 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_27 <= DFT_regdelays1_26; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_28 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_28 <= DFT_regdelays1_27; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_29 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_29 <= DFT_regdelays1_28; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_30 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_30 <= DFT_regdelays1_29; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_31 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_31 <= DFT_regdelays1_30; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_32 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_32 <= DFT_regdelays1_31; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_33 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_33 <= DFT_regdelays1_32; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_34 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_34 <= DFT_regdelays1_33; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_35 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_35 <= DFT_regdelays1_34; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6474:35]
      DFT_regdelays1_36 <= 1'h0; // @[FFTDesigns.scala 6474:35]
    end else begin
      DFT_regdelays1_36 <= DFT_regdelays1_35; // @[FFTDesigns.scala 6538:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6475:35]
      DFT_regdelays2_0 <= 1'h0; // @[FFTDesigns.scala 6475:35]
    end else begin
      DFT_regdelays2_0 <= Twid_regdelays_1; // @[FFTDesigns.scala 6544:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6475:35]
      DFT_regdelays2_1 <= 1'h0; // @[FFTDesigns.scala 6475:35]
    end else begin
      DFT_regdelays2_1 <= DFT_regdelays2_0; // @[FFTDesigns.scala 6551:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6475:35]
      DFT_regdelays2_2 <= 1'h0; // @[FFTDesigns.scala 6475:35]
    end else begin
      DFT_regdelays2_2 <= DFT_regdelays2_1; // @[FFTDesigns.scala 6551:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6475:35]
      DFT_regdelays2_3 <= 1'h0; // @[FFTDesigns.scala 6475:35]
    end else begin
      DFT_regdelays2_3 <= DFT_regdelays2_2; // @[FFTDesigns.scala 6551:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6476:35]
      Twid_regdelays_0 <= 1'h0; // @[FFTDesigns.scala 6476:35]
    end else begin
      Twid_regdelays_0 <= Perm_regdelays1_1_11; // @[FFTDesigns.scala 6523:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6476:35]
      Twid_regdelays_1 <= 1'h0; // @[FFTDesigns.scala 6476:35]
    end else begin
      Twid_regdelays_1 <= Twid_regdelays_0; // @[FFTDesigns.scala 6527:29]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_0 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_0 <= io_in_ready; // @[FFTDesigns.scala 6484:37]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_1 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_1 <= Perm_regdelays1_0_0; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_2 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_2 <= Perm_regdelays1_0_1; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_3 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_3 <= Perm_regdelays1_0_2; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_4 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_4 <= Perm_regdelays1_0_3; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_5 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_5 <= Perm_regdelays1_0_4; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_6 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_6 <= Perm_regdelays1_0_5; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_7 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_7 <= Perm_regdelays1_0_6; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_8 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_8 <= Perm_regdelays1_0_7; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_9 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_9 <= Perm_regdelays1_0_8; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_10 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_10 <= Perm_regdelays1_0_9; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_0_11 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_0_11 <= Perm_regdelays1_0_10; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_0 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_0 <= DFT_regdelays1_36; // @[FFTDesigns.scala 6488:37]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_1 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_1 <= Perm_regdelays1_1_0; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_2 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_2 <= Perm_regdelays1_1_1; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_3 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_3 <= Perm_regdelays1_1_2; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_4 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_4 <= Perm_regdelays1_1_3; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_5 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_5 <= Perm_regdelays1_1_4; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_6 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_6 <= Perm_regdelays1_1_5; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_7 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_7 <= Perm_regdelays1_1_6; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_8 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_8 <= Perm_regdelays1_1_7; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_9 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_9 <= Perm_regdelays1_1_8; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_10 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_10 <= Perm_regdelays1_1_9; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_1_11 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_1_11 <= Perm_regdelays1_1_10; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_0 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_0 <= DFT_regdelays2_3; // @[FFTDesigns.scala 6492:37]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_1 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_1 <= Perm_regdelays1_2_0; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_2 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_2 <= Perm_regdelays1_2_1; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_3 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_3 <= Perm_regdelays1_2_2; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_4 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_4 <= Perm_regdelays1_2_3; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_5 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_5 <= Perm_regdelays1_2_4; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_6 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_6 <= Perm_regdelays1_2_5; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_7 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_7 <= Perm_regdelays1_2_6; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_8 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_8 <= Perm_regdelays1_2_7; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_9 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_9 <= Perm_regdelays1_2_8; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_10 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_10 <= Perm_regdelays1_2_9; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6477:36]
      Perm_regdelays1_2_11 <= 1'h0; // @[FFTDesigns.scala 6477:36]
    end else begin
      Perm_regdelays1_2_11 <= Perm_regdelays1_2_10; // @[FFTDesigns.scala 6501:35]
    end
    if (reset) begin // @[FFTDesigns.scala 6478:33]
      out_regdelay <= 1'h0; // @[FFTDesigns.scala 6478:33]
    end else begin
      out_regdelay <= Perm_regdelays1_2_11; // @[FFTDesigns.scala 6554:20]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_0_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_0_Re <= PermutationsWithStreaming_mr_1_io_out_0_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_0_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_0_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_0_Im <= PermutationsWithStreaming_mr_1_io_out_0_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_0_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_1_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_1_Re <= PermutationsWithStreaming_mr_1_io_out_1_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_1_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_1_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_1_Im <= PermutationsWithStreaming_mr_1_io_out_1_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_1_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_2_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_2_Re <= PermutationsWithStreaming_mr_1_io_out_2_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_2_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_2_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_2_Im <= PermutationsWithStreaming_mr_1_io_out_2_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_2_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_3_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_3_Re <= PermutationsWithStreaming_mr_1_io_out_3_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_3_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_3_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_3_Im <= PermutationsWithStreaming_mr_1_io_out_3_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_3_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_4_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_4_Re <= PermutationsWithStreaming_mr_1_io_out_4_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_4_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_4_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_4_Im <= PermutationsWithStreaming_mr_1_io_out_4_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_4_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_5_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_5_Re <= PermutationsWithStreaming_mr_1_io_out_5_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_5_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_5_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_5_Im <= PermutationsWithStreaming_mr_1_io_out_5_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_5_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_6_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_6_Re <= PermutationsWithStreaming_mr_1_io_out_6_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_6_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_6_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_6_Im <= PermutationsWithStreaming_mr_1_io_out_6_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_6_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_7_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_7_Re <= PermutationsWithStreaming_mr_1_io_out_7_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_7_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_7_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_7_Im <= PermutationsWithStreaming_mr_1_io_out_7_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_7_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_8_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_8_Re <= PermutationsWithStreaming_mr_1_io_out_8_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_8_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_8_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_8_Im <= PermutationsWithStreaming_mr_1_io_out_8_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_8_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_9_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_9_Re <= PermutationsWithStreaming_mr_1_io_out_9_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_9_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_9_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_9_Im <= PermutationsWithStreaming_mr_1_io_out_9_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_9_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_10_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_10_Re <= PermutationsWithStreaming_mr_1_io_out_10_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_10_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_10_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_10_Im <= PermutationsWithStreaming_mr_1_io_out_10_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_10_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_11_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_11_Re <= PermutationsWithStreaming_mr_1_io_out_11_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_11_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_11_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_11_Im <= PermutationsWithStreaming_mr_1_io_out_11_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_11_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_12_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_12_Re <= PermutationsWithStreaming_mr_1_io_out_12_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_12_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_12_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_12_Im <= PermutationsWithStreaming_mr_1_io_out_12_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_12_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_13_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_13_Re <= PermutationsWithStreaming_mr_1_io_out_13_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_13_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_13_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_13_Im <= PermutationsWithStreaming_mr_1_io_out_13_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_13_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_14_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_14_Re <= PermutationsWithStreaming_mr_1_io_out_14_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_14_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_14_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_14_Im <= PermutationsWithStreaming_mr_1_io_out_14_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_14_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_15_Re <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_15_Re <= PermutationsWithStreaming_mr_1_io_out_15_Re; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_15_Re <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
    if (reset) begin // @[FFTDesigns.scala 6479:28]
      results_15_Im <= 32'h0; // @[FFTDesigns.scala 6479:28]
    end else if (Perm_regdelays1_2_11) begin // @[FFTDesigns.scala 6555:49]
      results_15_Im <= PermutationsWithStreaming_mr_1_io_out_15_Im; // @[FFTDesigns.scala 6556:17]
    end else begin
      results_15_Im <= 32'h0; // @[FFTDesigns.scala 6558:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DFT_regdelays1_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  DFT_regdelays1_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  DFT_regdelays1_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  DFT_regdelays1_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  DFT_regdelays1_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  DFT_regdelays1_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  DFT_regdelays1_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  DFT_regdelays1_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  DFT_regdelays1_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  DFT_regdelays1_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  DFT_regdelays1_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  DFT_regdelays1_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  DFT_regdelays1_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  DFT_regdelays1_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  DFT_regdelays1_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  DFT_regdelays1_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  DFT_regdelays1_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  DFT_regdelays1_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  DFT_regdelays1_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  DFT_regdelays1_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  DFT_regdelays1_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  DFT_regdelays1_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  DFT_regdelays1_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  DFT_regdelays1_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  DFT_regdelays1_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  DFT_regdelays1_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  DFT_regdelays1_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  DFT_regdelays1_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  DFT_regdelays1_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  DFT_regdelays1_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  DFT_regdelays1_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  DFT_regdelays1_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  DFT_regdelays1_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  DFT_regdelays1_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  DFT_regdelays1_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  DFT_regdelays1_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  DFT_regdelays1_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  DFT_regdelays2_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  DFT_regdelays2_1 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  DFT_regdelays2_2 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  DFT_regdelays2_3 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  Twid_regdelays_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  Twid_regdelays_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  Perm_regdelays1_0_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  Perm_regdelays1_0_1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  Perm_regdelays1_0_2 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  Perm_regdelays1_0_3 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  Perm_regdelays1_0_4 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  Perm_regdelays1_0_5 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  Perm_regdelays1_0_6 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  Perm_regdelays1_0_7 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  Perm_regdelays1_0_8 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  Perm_regdelays1_0_9 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  Perm_regdelays1_0_10 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  Perm_regdelays1_0_11 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  Perm_regdelays1_1_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  Perm_regdelays1_1_1 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  Perm_regdelays1_1_2 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  Perm_regdelays1_1_3 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  Perm_regdelays1_1_4 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  Perm_regdelays1_1_5 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  Perm_regdelays1_1_6 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  Perm_regdelays1_1_7 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  Perm_regdelays1_1_8 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  Perm_regdelays1_1_9 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  Perm_regdelays1_1_10 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  Perm_regdelays1_1_11 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  Perm_regdelays1_2_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  Perm_regdelays1_2_1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  Perm_regdelays1_2_2 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  Perm_regdelays1_2_3 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  Perm_regdelays1_2_4 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  Perm_regdelays1_2_5 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  Perm_regdelays1_2_6 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  Perm_regdelays1_2_7 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  Perm_regdelays1_2_8 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  Perm_regdelays1_2_9 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  Perm_regdelays1_2_10 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  Perm_regdelays1_2_11 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  out_regdelay = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  results_0_Re = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  results_0_Im = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  results_1_Re = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  results_1_Im = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  results_2_Re = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  results_2_Im = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  results_3_Re = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  results_3_Im = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  results_4_Re = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  results_4_Im = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  results_5_Re = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  results_5_Im = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  results_6_Re = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  results_6_Im = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  results_7_Re = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  results_7_Im = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  results_8_Re = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  results_8_Im = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  results_9_Re = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  results_9_Im = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  results_10_Re = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  results_10_Im = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  results_11_Re = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  results_11_Im = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  results_12_Re = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  results_12_Im = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  results_13_Re = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  results_13_Im = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  results_14_Re = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  results_14_Im = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  results_15_Re = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  results_15_Im = _RAND_111[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

